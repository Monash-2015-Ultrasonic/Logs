// NIOS_SYSTEMV3.v

// Generated using ACDS version 13.0sp1 232 at 2015.10.23.09:54:52

`timescale 1 ps / 1 ps
module NIOS_SYSTEMV3 (
		input  wire        clk_clk,                                           //                   clk.clk
		input  wire        reset_reset_n,                                     //                 reset.reset_n
		output wire        lcd_RS,                                            //                   lcd.RS
		output wire        lcd_RW,                                            //                      .RW
		inout  wire [7:0]  lcd_data,                                          //                      .data
		output wire        lcd_E,                                             //                      .E
		output wire        adc_on_export,                                     //                adc_on.export
		output wire [15:0] fifo_adc_data_export,                              //         fifo_adc_data.export
		output wire        fifo_adc_data_valid_export,                        //   fifo_adc_data_valid.export
		output wire        fifo_rst_export,                                   //              fifo_rst.export
		output wire        subtractor_on_export,                              //         subtractor_on.export
		output wire        ch0_timer_rst_export,                              //         ch0_timer_rst.export
		output wire        detector_on_export,                                //           detector_on.export
		input  wire        menu_export,                                       //                  menu.export
		input  wire        menu_up_export,                                    //               menu_up.export
		input  wire        menu_down_export,                                  //             menu_down.export
		output wire [23:0] ch0_thresh_export,                                 //            ch0_thresh.export
		output wire        ch0_rd_peak_export,                                //           ch0_rd_peak.export
		input  wire        ch0_peak_found_export,                             //        ch0_peak_found.export
		input  wire [13:0] ch0_yn1_u_export,                                  //             ch0_yn1_u.export
		input  wire [31:0] ch0_yn1_mu_export,                                 //            ch0_yn1_mu.export
		input  wire [31:0] ch0_yn1_ml_export,                                 //            ch0_yn1_ml.export
		input  wire [31:0] ch0_yn1_l_export,                                  //             ch0_yn1_l.export
		input  wire [13:0] ch0_time_export,                                   //              ch0_time.export
		input  wire [31:0] ch0_yn2_l_export,                                  //             ch0_yn2_l.export
		input  wire [31:0] ch0_yn2_ml_export,                                 //            ch0_yn2_ml.export
		input  wire [31:0] ch0_yn2_mu_export,                                 //            ch0_yn2_mu.export
		input  wire [13:0] ch0_yn2_u_export,                                  //             ch0_yn2_u.export
		input  wire [13:0] ch0_yn3_u_export,                                  //             ch0_yn3_u.export
		input  wire [31:0] ch0_yn3_mu_export,                                 //            ch0_yn3_mu.export
		input  wire [31:0] ch0_yn3_ml_export,                                 //            ch0_yn3_ml.export
		input  wire [31:0] ch0_yn3_l_export,                                  //             ch0_yn3_l.export
		output wire        ch1_timer_rst_export,                              //         ch1_timer_rst.export
		output wire [23:0] ch1_thresh_export,                                 //            ch1_thresh.export
		output wire        ch1_rd_peak_export,                                //           ch1_rd_peak.export
		input  wire        ch1_peak_found_export,                             //        ch1_peak_found.export
		input  wire [13:0] ch1_time_export,                                   //              ch1_time.export
		input  wire [13:0] ch1_yn1_u_export,                                  //             ch1_yn1_u.export
		input  wire [31:0] ch1_yn1_mu_export,                                 //            ch1_yn1_mu.export
		input  wire [31:0] ch1_yn1_ml_export,                                 //            ch1_yn1_ml.export
		input  wire [31:0] ch1_yn1_l_export,                                  //             ch1_yn1_l.export
		input  wire [13:0] ch1_yn2_u_export,                                  //             ch1_yn2_u.export
		input  wire [31:0] ch1_yn2_mu_export,                                 //            ch1_yn2_mu.export
		input  wire [31:0] ch1_yn2_ml_export,                                 //            ch1_yn2_ml.export
		input  wire [31:0] ch1_yn2_l_export,                                  //             ch1_yn2_l.export
		input  wire [13:0] ch1_yn3_u_export,                                  //             ch1_yn3_u.export
		input  wire [31:0] ch1_yn3_mu_export,                                 //            ch1_yn3_mu.export
		input  wire [31:0] ch1_yn3_ml_export,                                 //            ch1_yn3_ml.export
		input  wire [31:0] ch1_yn3_l_export,                                  //             ch1_yn3_l.export
		output wire        ch2_timer_rst_export,                              //         ch2_timer_rst.export
		output wire [23:0] ch2_thresh_export,                                 //            ch2_thresh.export
		output wire        ch2_rd_peak_export,                                //           ch2_rd_peak.export
		input  wire        ch2_peak_found_export,                             //        ch2_peak_found.export
		input  wire [13:0] ch2_time_export,                                   //              ch2_time.export
		input  wire [13:0] ch2_yn1_u_export,                                  //             ch2_yn1_u.export
		input  wire [31:0] ch2_yn1_mu_export,                                 //            ch2_yn1_mu.export
		input  wire [31:0] ch2_yn1_ml_export,                                 //            ch2_yn1_ml.export
		input  wire [31:0] ch2_yn1_l_export,                                  //             ch2_yn1_l.export
		input  wire [13:0] ch2_yn2_u_export,                                  //             ch2_yn2_u.export
		input  wire [31:0] ch2_yn2_mu_export,                                 //            ch2_yn2_mu.export
		input  wire [31:0] ch2_yn2_ml_export,                                 //            ch2_yn2_ml.export
		input  wire [31:0] ch2_yn2_l_export,                                  //             ch2_yn2_l.export
		input  wire [13:0] ch2_yn3_u_export,                                  //             ch2_yn3_u.export
		input  wire [31:0] ch2_yn3_mu_export,                                 //            ch2_yn3_mu.export
		input  wire [31:0] ch2_yn3_ml_export,                                 //            ch2_yn3_ml.export
		input  wire [31:0] ch2_yn3_l_export,                                  //             ch2_yn3_l.export
		input  wire [31:0] ch3_yn3_l_export,                                  //             ch3_yn3_l.export
		input  wire [31:0] ch3_yn3_ml_export,                                 //            ch3_yn3_ml.export
		input  wire [31:0] ch3_yn3_mu_export,                                 //            ch3_yn3_mu.export
		input  wire [13:0] ch3_yn3_u_export,                                  //             ch3_yn3_u.export
		input  wire [31:0] ch3_yn2_l_export,                                  //             ch3_yn2_l.export
		input  wire [31:0] ch3_yn2_ml_export,                                 //            ch3_yn2_ml.export
		input  wire [31:0] ch3_yn2_mu_export,                                 //            ch3_yn2_mu.export
		input  wire [13:0] ch3_yn2_u_export,                                  //             ch3_yn2_u.export
		input  wire [31:0] ch3_yn1_l_export,                                  //             ch3_yn1_l.export
		input  wire [31:0] ch3_yn1_ml_export,                                 //            ch3_yn1_ml.export
		input  wire [31:0] ch3_yn1_mu_export,                                 //            ch3_yn1_mu.export
		input  wire [13:0] ch3_yn1_u_export,                                  //             ch3_yn1_u.export
		input  wire [13:0] ch3_time_export,                                   //              ch3_time.export
		output wire        ch3_timer_rst_export,                              //         ch3_timer_rst.export
		output wire [23:0] ch3_thresh_export,                                 //            ch3_thresh.export
		output wire        ch3_rd_peak_export,                                //           ch3_rd_peak.export
		input  wire        ch3_peak_found_export,                             //        ch3_peak_found.export
		input  wire [31:0] ch4_yn3_l_export,                                  //             ch4_yn3_l.export
		input  wire [31:0] ch4_yn3_ml_export,                                 //            ch4_yn3_ml.export
		input  wire [31:0] ch4_yn3_mu_export,                                 //            ch4_yn3_mu.export
		input  wire [13:0] ch4_yn3_u_export,                                  //             ch4_yn3_u.export
		input  wire [31:0] ch4_yn2_l_export,                                  //             ch4_yn2_l.export
		input  wire [31:0] ch4_yn2_ml_export,                                 //            ch4_yn2_ml.export
		input  wire [31:0] ch4_yn2_mu_export,                                 //            ch4_yn2_mu.export
		input  wire [13:0] ch4_yn2_u_export,                                  //             ch4_yn2_u.export
		input  wire [31:0] ch4_yn1_l_export,                                  //             ch4_yn1_l.export
		input  wire [31:0] ch4_yn1_ml_export,                                 //            ch4_yn1_ml.export
		input  wire [31:0] ch4_yn1_mu_export,                                 //            ch4_yn1_mu.export
		input  wire [13:0] ch4_yn1_u_export,                                  //             ch4_yn1_u.export
		input  wire [13:0] ch4_time_export,                                   //              ch4_time.export
		input  wire        ch4_peak_found_export,                             //        ch4_peak_found.export
		output wire        ch4_timer_rst_export,                              //         ch4_timer_rst.export
		output wire [23:0] ch4_thresh_export,                                 //            ch4_thresh.export
		output wire        ch4_rd_peak_export,                                //           ch4_rd_peak.export
		output wire [0:0]  tristate_bridge_ssram_bwe_n_to_the_ssram,          // tristate_bridge_ssram.bwe_n_to_the_ssram
		output wire [0:0]  tristate_bridge_ssram_reset_n_to_the_ssram,        //                      .reset_n_to_the_ssram
		output wire [0:0]  tristate_bridge_ssram_chipenable1_n_to_the_ssram,  //                      .chipenable1_n_to_the_ssram
		output wire [3:0]  tristate_bridge_ssram_bw_n_to_the_ssram,           //                      .bw_n_to_the_ssram
		output wire [0:0]  tristate_bridge_ssram_outputenable_n_to_the_ssram, //                      .outputenable_n_to_the_ssram
		output wire [0:0]  tristate_bridge_ssram_adsc_n_to_the_ssram,         //                      .adsc_n_to_the_ssram
		output wire [20:0] tristate_bridge_ssram_address_to_the_ssram,        //                      .address_to_the_ssram
		inout  wire [31:0] tristate_bridge_ssram_data_to_and_from_the_ssram   //                      .data_to_and_from_the_ssram
	);

	wire          nios_cpu_jtag_debug_module_reset_reset;                                                           // NIOS_CPU:jtag_debug_module_resetrequest -> [CH2_YN1_L:reset_n, CH2_YN1_L_s1_translator:reset, CH2_YN1_L_s1_translator_avalon_universal_slave_0_agent:reset, CH2_YN1_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, id_router_056:reset, rsp_xbar_demux_056:reset, rst_controller_001:reset_in0]
	wire          tristate_bridge_ssram_pinsharer_tcm_data_to_and_from_the_ssram_outen;                             // tristate_bridge_ssram_pinSharer:data_to_and_from_the_ssram_outen -> tristate_bridge_ssram:tcs_data_to_and_from_the_ssram_outen
	wire    [0:0] tristate_bridge_ssram_pinsharer_tcm_outputenable_n_to_the_ssram_out;                              // tristate_bridge_ssram_pinSharer:outputenable_n_to_the_ssram -> tristate_bridge_ssram:tcs_outputenable_n_to_the_ssram
	wire          tristate_bridge_ssram_pinsharer_tcm_grant;                                                        // tristate_bridge_ssram:grant -> tristate_bridge_ssram_pinSharer:grant
	wire          tristate_bridge_ssram_pinsharer_tcm_request;                                                      // tristate_bridge_ssram_pinSharer:request -> tristate_bridge_ssram:request
	wire   [31:0] tristate_bridge_ssram_pinsharer_tcm_data_to_and_from_the_ssram_in;                                // tristate_bridge_ssram:tcs_data_to_and_from_the_ssram_in -> tristate_bridge_ssram_pinSharer:data_to_and_from_the_ssram_in
	wire   [31:0] tristate_bridge_ssram_pinsharer_tcm_data_to_and_from_the_ssram_out;                               // tristate_bridge_ssram_pinSharer:data_to_and_from_the_ssram -> tristate_bridge_ssram:tcs_data_to_and_from_the_ssram
	wire    [0:0] tristate_bridge_ssram_pinsharer_tcm_bwe_n_to_the_ssram_out;                                       // tristate_bridge_ssram_pinSharer:bwe_n_to_the_ssram -> tristate_bridge_ssram:tcs_bwe_n_to_the_ssram
	wire    [0:0] tristate_bridge_ssram_pinsharer_tcm_adsc_n_to_the_ssram_out;                                      // tristate_bridge_ssram_pinSharer:adsc_n_to_the_ssram -> tristate_bridge_ssram:tcs_adsc_n_to_the_ssram
	wire    [0:0] tristate_bridge_ssram_pinsharer_tcm_reset_n_to_the_ssram_out;                                     // tristate_bridge_ssram_pinSharer:reset_n_to_the_ssram -> tristate_bridge_ssram:tcs_reset_n_to_the_ssram
	wire    [0:0] tristate_bridge_ssram_pinsharer_tcm_chipenable1_n_to_the_ssram_out;                               // tristate_bridge_ssram_pinSharer:chipenable1_n_to_the_ssram -> tristate_bridge_ssram:tcs_chipenable1_n_to_the_ssram
	wire   [20:0] tristate_bridge_ssram_pinsharer_tcm_address_to_the_ssram_out;                                     // tristate_bridge_ssram_pinSharer:address_to_the_ssram -> tristate_bridge_ssram:tcs_address_to_the_ssram
	wire    [3:0] tristate_bridge_ssram_pinsharer_tcm_bw_n_to_the_ssram_out;                                        // tristate_bridge_ssram_pinSharer:bw_n_to_the_ssram -> tristate_bridge_ssram:tcs_bw_n_to_the_ssram
	wire          ssram_tcm_chipselect_n_out;                                                                       // SSRAM:tcm_chipselect_n_out -> tristate_bridge_ssram_pinSharer:tcs0_chipselect_n_out
	wire          ssram_tcm_grant;                                                                                  // tristate_bridge_ssram_pinSharer:tcs0_grant -> SSRAM:tcm_grant
	wire          ssram_tcm_data_outen;                                                                             // SSRAM:tcm_data_outen -> tristate_bridge_ssram_pinSharer:tcs0_data_outen
	wire          ssram_tcm_reset_n_out;                                                                            // SSRAM:tcm_reset_n_out -> tristate_bridge_ssram_pinSharer:tcs0_reset_n_out
	wire          ssram_tcm_outputenable_n_out;                                                                     // SSRAM:tcm_outputenable_n_out -> tristate_bridge_ssram_pinSharer:tcs0_outputenable_n_out
	wire          ssram_tcm_request;                                                                                // SSRAM:tcm_request -> tristate_bridge_ssram_pinSharer:tcs0_request
	wire   [31:0] ssram_tcm_data_out;                                                                               // SSRAM:tcm_data_out -> tristate_bridge_ssram_pinSharer:tcs0_data_out
	wire          ssram_tcm_write_n_out;                                                                            // SSRAM:tcm_write_n_out -> tristate_bridge_ssram_pinSharer:tcs0_write_n_out
	wire   [20:0] ssram_tcm_address_out;                                                                            // SSRAM:tcm_address_out -> tristate_bridge_ssram_pinSharer:tcs0_address_out
	wire   [31:0] ssram_tcm_data_in;                                                                                // tristate_bridge_ssram_pinSharer:tcs0_data_in -> SSRAM:tcm_data_in
	wire          ssram_tcm_begintransfer_n_out;                                                                    // SSRAM:tcm_begintransfer_n_out -> tristate_bridge_ssram_pinSharer:tcs0_begintransfer_n_out
	wire    [3:0] ssram_tcm_byteenable_n_out;                                                                       // SSRAM:tcm_byteenable_n_out -> tristate_bridge_ssram_pinSharer:tcs0_byteenable_n_out
	wire          nios_cpu_instruction_master_waitrequest;                                                          // NIOS_CPU_instruction_master_translator:av_waitrequest -> NIOS_CPU:i_waitrequest
	wire   [21:0] nios_cpu_instruction_master_address;                                                              // NIOS_CPU:i_address -> NIOS_CPU_instruction_master_translator:av_address
	wire          nios_cpu_instruction_master_read;                                                                 // NIOS_CPU:i_read -> NIOS_CPU_instruction_master_translator:av_read
	wire   [31:0] nios_cpu_instruction_master_readdata;                                                             // NIOS_CPU_instruction_master_translator:av_readdata -> NIOS_CPU:i_readdata
	wire          nios_cpu_data_master_waitrequest;                                                                 // NIOS_CPU_data_master_translator:av_waitrequest -> NIOS_CPU:d_waitrequest
	wire   [31:0] nios_cpu_data_master_writedata;                                                                   // NIOS_CPU:d_writedata -> NIOS_CPU_data_master_translator:av_writedata
	wire   [21:0] nios_cpu_data_master_address;                                                                     // NIOS_CPU:d_address -> NIOS_CPU_data_master_translator:av_address
	wire          nios_cpu_data_master_write;                                                                       // NIOS_CPU:d_write -> NIOS_CPU_data_master_translator:av_write
	wire          nios_cpu_data_master_read;                                                                        // NIOS_CPU:d_read -> NIOS_CPU_data_master_translator:av_read
	wire   [31:0] nios_cpu_data_master_readdata;                                                                    // NIOS_CPU_data_master_translator:av_readdata -> NIOS_CPU:d_readdata
	wire          nios_cpu_data_master_debugaccess;                                                                 // NIOS_CPU:jtag_debug_module_debugaccess_to_roms -> NIOS_CPU_data_master_translator:av_debugaccess
	wire    [3:0] nios_cpu_data_master_byteenable;                                                                  // NIOS_CPU:d_byteenable -> NIOS_CPU_data_master_translator:av_byteenable
	wire          nios_cpu_jtag_debug_module_translator_avalon_anti_slave_0_waitrequest;                            // NIOS_CPU:jtag_debug_module_waitrequest -> NIOS_CPU_jtag_debug_module_translator:av_waitrequest
	wire   [31:0] nios_cpu_jtag_debug_module_translator_avalon_anti_slave_0_writedata;                              // NIOS_CPU_jtag_debug_module_translator:av_writedata -> NIOS_CPU:jtag_debug_module_writedata
	wire    [8:0] nios_cpu_jtag_debug_module_translator_avalon_anti_slave_0_address;                                // NIOS_CPU_jtag_debug_module_translator:av_address -> NIOS_CPU:jtag_debug_module_address
	wire          nios_cpu_jtag_debug_module_translator_avalon_anti_slave_0_write;                                  // NIOS_CPU_jtag_debug_module_translator:av_write -> NIOS_CPU:jtag_debug_module_write
	wire          nios_cpu_jtag_debug_module_translator_avalon_anti_slave_0_read;                                   // NIOS_CPU_jtag_debug_module_translator:av_read -> NIOS_CPU:jtag_debug_module_read
	wire   [31:0] nios_cpu_jtag_debug_module_translator_avalon_anti_slave_0_readdata;                               // NIOS_CPU:jtag_debug_module_readdata -> NIOS_CPU_jtag_debug_module_translator:av_readdata
	wire          nios_cpu_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess;                            // NIOS_CPU_jtag_debug_module_translator:av_debugaccess -> NIOS_CPU:jtag_debug_module_debugaccess
	wire    [3:0] nios_cpu_jtag_debug_module_translator_avalon_anti_slave_0_byteenable;                             // NIOS_CPU_jtag_debug_module_translator:av_byteenable -> NIOS_CPU:jtag_debug_module_byteenable
	wire   [31:0] ram_s1_translator_avalon_anti_slave_0_writedata;                                                  // RAM_s1_translator:av_writedata -> RAM:writedata
	wire   [10:0] ram_s1_translator_avalon_anti_slave_0_address;                                                    // RAM_s1_translator:av_address -> RAM:address
	wire          ram_s1_translator_avalon_anti_slave_0_chipselect;                                                 // RAM_s1_translator:av_chipselect -> RAM:chipselect
	wire          ram_s1_translator_avalon_anti_slave_0_clken;                                                      // RAM_s1_translator:av_clken -> RAM:clken
	wire          ram_s1_translator_avalon_anti_slave_0_write;                                                      // RAM_s1_translator:av_write -> RAM:write
	wire   [31:0] ram_s1_translator_avalon_anti_slave_0_readdata;                                                   // RAM:readdata -> RAM_s1_translator:av_readdata
	wire    [3:0] ram_s1_translator_avalon_anti_slave_0_byteenable;                                                 // RAM_s1_translator:av_byteenable -> RAM:byteenable
	wire          ssram_uas_translator_avalon_anti_slave_0_waitrequest;                                             // SSRAM:uas_waitrequest -> SSRAM_uas_translator:av_waitrequest
	wire    [2:0] ssram_uas_translator_avalon_anti_slave_0_burstcount;                                              // SSRAM_uas_translator:av_burstcount -> SSRAM:uas_burstcount
	wire   [31:0] ssram_uas_translator_avalon_anti_slave_0_writedata;                                               // SSRAM_uas_translator:av_writedata -> SSRAM:uas_writedata
	wire   [20:0] ssram_uas_translator_avalon_anti_slave_0_address;                                                 // SSRAM_uas_translator:av_address -> SSRAM:uas_address
	wire          ssram_uas_translator_avalon_anti_slave_0_lock;                                                    // SSRAM_uas_translator:av_lock -> SSRAM:uas_lock
	wire          ssram_uas_translator_avalon_anti_slave_0_write;                                                   // SSRAM_uas_translator:av_write -> SSRAM:uas_write
	wire          ssram_uas_translator_avalon_anti_slave_0_read;                                                    // SSRAM_uas_translator:av_read -> SSRAM:uas_read
	wire   [31:0] ssram_uas_translator_avalon_anti_slave_0_readdata;                                                // SSRAM:uas_readdata -> SSRAM_uas_translator:av_readdata
	wire          ssram_uas_translator_avalon_anti_slave_0_debugaccess;                                             // SSRAM_uas_translator:av_debugaccess -> SSRAM:uas_debugaccess
	wire          ssram_uas_translator_avalon_anti_slave_0_readdatavalid;                                           // SSRAM:uas_readdatavalid -> SSRAM_uas_translator:av_readdatavalid
	wire    [3:0] ssram_uas_translator_avalon_anti_slave_0_byteenable;                                              // SSRAM_uas_translator:av_byteenable -> SSRAM:uas_byteenable
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest;                           // JTAG_UART:av_waitrequest -> JTAG_UART_avalon_jtag_slave_translator:av_waitrequest
	wire   [31:0] jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata;                             // JTAG_UART_avalon_jtag_slave_translator:av_writedata -> JTAG_UART:av_writedata
	wire    [0:0] jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_address;                               // JTAG_UART_avalon_jtag_slave_translator:av_address -> JTAG_UART:av_address
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect;                            // JTAG_UART_avalon_jtag_slave_translator:av_chipselect -> JTAG_UART:av_chipselect
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_write;                                 // JTAG_UART_avalon_jtag_slave_translator:av_write -> JTAG_UART:av_write_n
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_read;                                  // JTAG_UART_avalon_jtag_slave_translator:av_read -> JTAG_UART:av_read_n
	wire   [31:0] jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata;                              // JTAG_UART:av_readdata -> JTAG_UART_avalon_jtag_slave_translator:av_readdata
	wire    [7:0] lcd_control_slave_translator_avalon_anti_slave_0_writedata;                                       // LCD_control_slave_translator:av_writedata -> LCD:writedata
	wire    [1:0] lcd_control_slave_translator_avalon_anti_slave_0_address;                                         // LCD_control_slave_translator:av_address -> LCD:address
	wire          lcd_control_slave_translator_avalon_anti_slave_0_write;                                           // LCD_control_slave_translator:av_write -> LCD:write
	wire          lcd_control_slave_translator_avalon_anti_slave_0_read;                                            // LCD_control_slave_translator:av_read -> LCD:read
	wire    [7:0] lcd_control_slave_translator_avalon_anti_slave_0_readdata;                                        // LCD:readdata -> LCD_control_slave_translator:av_readdata
	wire          lcd_control_slave_translator_avalon_anti_slave_0_begintransfer;                                   // LCD_control_slave_translator:av_begintransfer -> LCD:begintransfer
	wire   [31:0] adc_on_s1_translator_avalon_anti_slave_0_writedata;                                               // ADC_ON_s1_translator:av_writedata -> ADC_ON:writedata
	wire    [1:0] adc_on_s1_translator_avalon_anti_slave_0_address;                                                 // ADC_ON_s1_translator:av_address -> ADC_ON:address
	wire          adc_on_s1_translator_avalon_anti_slave_0_chipselect;                                              // ADC_ON_s1_translator:av_chipselect -> ADC_ON:chipselect
	wire          adc_on_s1_translator_avalon_anti_slave_0_write;                                                   // ADC_ON_s1_translator:av_write -> ADC_ON:write_n
	wire   [31:0] adc_on_s1_translator_avalon_anti_slave_0_readdata;                                                // ADC_ON:readdata -> ADC_ON_s1_translator:av_readdata
	wire   [31:0] fifo_adc_data_s1_translator_avalon_anti_slave_0_writedata;                                        // FIFO_ADC_DATA_s1_translator:av_writedata -> FIFO_ADC_DATA:writedata
	wire    [1:0] fifo_adc_data_s1_translator_avalon_anti_slave_0_address;                                          // FIFO_ADC_DATA_s1_translator:av_address -> FIFO_ADC_DATA:address
	wire          fifo_adc_data_s1_translator_avalon_anti_slave_0_chipselect;                                       // FIFO_ADC_DATA_s1_translator:av_chipselect -> FIFO_ADC_DATA:chipselect
	wire          fifo_adc_data_s1_translator_avalon_anti_slave_0_write;                                            // FIFO_ADC_DATA_s1_translator:av_write -> FIFO_ADC_DATA:write_n
	wire   [31:0] fifo_adc_data_s1_translator_avalon_anti_slave_0_readdata;                                         // FIFO_ADC_DATA:readdata -> FIFO_ADC_DATA_s1_translator:av_readdata
	wire   [31:0] fifo_adc_data_valid_s1_translator_avalon_anti_slave_0_writedata;                                  // FIFO_ADC_DATA_VALID_s1_translator:av_writedata -> FIFO_ADC_DATA_VALID:writedata
	wire    [1:0] fifo_adc_data_valid_s1_translator_avalon_anti_slave_0_address;                                    // FIFO_ADC_DATA_VALID_s1_translator:av_address -> FIFO_ADC_DATA_VALID:address
	wire          fifo_adc_data_valid_s1_translator_avalon_anti_slave_0_chipselect;                                 // FIFO_ADC_DATA_VALID_s1_translator:av_chipselect -> FIFO_ADC_DATA_VALID:chipselect
	wire          fifo_adc_data_valid_s1_translator_avalon_anti_slave_0_write;                                      // FIFO_ADC_DATA_VALID_s1_translator:av_write -> FIFO_ADC_DATA_VALID:write_n
	wire   [31:0] fifo_adc_data_valid_s1_translator_avalon_anti_slave_0_readdata;                                   // FIFO_ADC_DATA_VALID:readdata -> FIFO_ADC_DATA_VALID_s1_translator:av_readdata
	wire   [31:0] fifo_rst_s1_translator_avalon_anti_slave_0_writedata;                                             // FIFO_RST_s1_translator:av_writedata -> FIFO_RST:writedata
	wire    [1:0] fifo_rst_s1_translator_avalon_anti_slave_0_address;                                               // FIFO_RST_s1_translator:av_address -> FIFO_RST:address
	wire          fifo_rst_s1_translator_avalon_anti_slave_0_chipselect;                                            // FIFO_RST_s1_translator:av_chipselect -> FIFO_RST:chipselect
	wire          fifo_rst_s1_translator_avalon_anti_slave_0_write;                                                 // FIFO_RST_s1_translator:av_write -> FIFO_RST:write_n
	wire   [31:0] fifo_rst_s1_translator_avalon_anti_slave_0_readdata;                                              // FIFO_RST:readdata -> FIFO_RST_s1_translator:av_readdata
	wire   [31:0] subtractor_on_s1_translator_avalon_anti_slave_0_writedata;                                        // SUBTRACTOR_ON_s1_translator:av_writedata -> SUBTRACTOR_ON:writedata
	wire    [1:0] subtractor_on_s1_translator_avalon_anti_slave_0_address;                                          // SUBTRACTOR_ON_s1_translator:av_address -> SUBTRACTOR_ON:address
	wire          subtractor_on_s1_translator_avalon_anti_slave_0_chipselect;                                       // SUBTRACTOR_ON_s1_translator:av_chipselect -> SUBTRACTOR_ON:chipselect
	wire          subtractor_on_s1_translator_avalon_anti_slave_0_write;                                            // SUBTRACTOR_ON_s1_translator:av_write -> SUBTRACTOR_ON:write_n
	wire   [31:0] subtractor_on_s1_translator_avalon_anti_slave_0_readdata;                                         // SUBTRACTOR_ON:readdata -> SUBTRACTOR_ON_s1_translator:av_readdata
	wire   [31:0] ch0_timer_rst_s1_translator_avalon_anti_slave_0_writedata;                                        // CH0_TIMER_RST_s1_translator:av_writedata -> CH0_TIMER_RST:writedata
	wire    [1:0] ch0_timer_rst_s1_translator_avalon_anti_slave_0_address;                                          // CH0_TIMER_RST_s1_translator:av_address -> CH0_TIMER_RST:address
	wire          ch0_timer_rst_s1_translator_avalon_anti_slave_0_chipselect;                                       // CH0_TIMER_RST_s1_translator:av_chipselect -> CH0_TIMER_RST:chipselect
	wire          ch0_timer_rst_s1_translator_avalon_anti_slave_0_write;                                            // CH0_TIMER_RST_s1_translator:av_write -> CH0_TIMER_RST:write_n
	wire   [31:0] ch0_timer_rst_s1_translator_avalon_anti_slave_0_readdata;                                         // CH0_TIMER_RST:readdata -> CH0_TIMER_RST_s1_translator:av_readdata
	wire   [31:0] detector_on_s1_translator_avalon_anti_slave_0_writedata;                                          // DETECTOR_ON_s1_translator:av_writedata -> DETECTOR_ON:writedata
	wire    [1:0] detector_on_s1_translator_avalon_anti_slave_0_address;                                            // DETECTOR_ON_s1_translator:av_address -> DETECTOR_ON:address
	wire          detector_on_s1_translator_avalon_anti_slave_0_chipselect;                                         // DETECTOR_ON_s1_translator:av_chipselect -> DETECTOR_ON:chipselect
	wire          detector_on_s1_translator_avalon_anti_slave_0_write;                                              // DETECTOR_ON_s1_translator:av_write -> DETECTOR_ON:write_n
	wire   [31:0] detector_on_s1_translator_avalon_anti_slave_0_readdata;                                           // DETECTOR_ON:readdata -> DETECTOR_ON_s1_translator:av_readdata
	wire    [1:0] menu_down_s1_translator_avalon_anti_slave_0_address;                                              // MENU_DOWN_s1_translator:av_address -> MENU_DOWN:address
	wire   [31:0] menu_down_s1_translator_avalon_anti_slave_0_readdata;                                             // MENU_DOWN:readdata -> MENU_DOWN_s1_translator:av_readdata
	wire   [31:0] menu_up_s1_translator_avalon_anti_slave_0_writedata;                                              // MENU_UP_s1_translator:av_writedata -> MENU_UP:writedata
	wire    [1:0] menu_up_s1_translator_avalon_anti_slave_0_address;                                                // MENU_UP_s1_translator:av_address -> MENU_UP:address
	wire          menu_up_s1_translator_avalon_anti_slave_0_chipselect;                                             // MENU_UP_s1_translator:av_chipselect -> MENU_UP:chipselect
	wire          menu_up_s1_translator_avalon_anti_slave_0_write;                                                  // MENU_UP_s1_translator:av_write -> MENU_UP:write_n
	wire   [31:0] menu_up_s1_translator_avalon_anti_slave_0_readdata;                                               // MENU_UP:readdata -> MENU_UP_s1_translator:av_readdata
	wire   [31:0] menu_s1_translator_avalon_anti_slave_0_writedata;                                                 // MENU_s1_translator:av_writedata -> MENU:writedata
	wire    [1:0] menu_s1_translator_avalon_anti_slave_0_address;                                                   // MENU_s1_translator:av_address -> MENU:address
	wire          menu_s1_translator_avalon_anti_slave_0_chipselect;                                                // MENU_s1_translator:av_chipselect -> MENU:chipselect
	wire          menu_s1_translator_avalon_anti_slave_0_write;                                                     // MENU_s1_translator:av_write -> MENU:write_n
	wire   [31:0] menu_s1_translator_avalon_anti_slave_0_readdata;                                                  // MENU:readdata -> MENU_s1_translator:av_readdata
	wire   [31:0] ch0_thresh_s1_translator_avalon_anti_slave_0_writedata;                                           // CH0_THRESH_s1_translator:av_writedata -> CH0_THRESH:writedata
	wire    [1:0] ch0_thresh_s1_translator_avalon_anti_slave_0_address;                                             // CH0_THRESH_s1_translator:av_address -> CH0_THRESH:address
	wire          ch0_thresh_s1_translator_avalon_anti_slave_0_chipselect;                                          // CH0_THRESH_s1_translator:av_chipselect -> CH0_THRESH:chipselect
	wire          ch0_thresh_s1_translator_avalon_anti_slave_0_write;                                               // CH0_THRESH_s1_translator:av_write -> CH0_THRESH:write_n
	wire   [31:0] ch0_thresh_s1_translator_avalon_anti_slave_0_readdata;                                            // CH0_THRESH:readdata -> CH0_THRESH_s1_translator:av_readdata
	wire   [31:0] ch0_rd_peak_s1_translator_avalon_anti_slave_0_writedata;                                          // CH0_RD_PEAK_s1_translator:av_writedata -> CH0_RD_PEAK:writedata
	wire    [1:0] ch0_rd_peak_s1_translator_avalon_anti_slave_0_address;                                            // CH0_RD_PEAK_s1_translator:av_address -> CH0_RD_PEAK:address
	wire          ch0_rd_peak_s1_translator_avalon_anti_slave_0_chipselect;                                         // CH0_RD_PEAK_s1_translator:av_chipselect -> CH0_RD_PEAK:chipselect
	wire          ch0_rd_peak_s1_translator_avalon_anti_slave_0_write;                                              // CH0_RD_PEAK_s1_translator:av_write -> CH0_RD_PEAK:write_n
	wire   [31:0] ch0_rd_peak_s1_translator_avalon_anti_slave_0_readdata;                                           // CH0_RD_PEAK:readdata -> CH0_RD_PEAK_s1_translator:av_readdata
	wire   [31:0] ch0_peak_found_s1_translator_avalon_anti_slave_0_writedata;                                       // CH0_PEAK_FOUND_s1_translator:av_writedata -> CH0_PEAK_FOUND:writedata
	wire    [1:0] ch0_peak_found_s1_translator_avalon_anti_slave_0_address;                                         // CH0_PEAK_FOUND_s1_translator:av_address -> CH0_PEAK_FOUND:address
	wire          ch0_peak_found_s1_translator_avalon_anti_slave_0_chipselect;                                      // CH0_PEAK_FOUND_s1_translator:av_chipselect -> CH0_PEAK_FOUND:chipselect
	wire          ch0_peak_found_s1_translator_avalon_anti_slave_0_write;                                           // CH0_PEAK_FOUND_s1_translator:av_write -> CH0_PEAK_FOUND:write_n
	wire   [31:0] ch0_peak_found_s1_translator_avalon_anti_slave_0_readdata;                                        // CH0_PEAK_FOUND:readdata -> CH0_PEAK_FOUND_s1_translator:av_readdata
	wire   [31:0] ch0_yn1_l_s1_translator_avalon_anti_slave_0_writedata;                                            // CH0_YN1_L_s1_translator:av_writedata -> CH0_YN1_L:writedata
	wire    [1:0] ch0_yn1_l_s1_translator_avalon_anti_slave_0_address;                                              // CH0_YN1_L_s1_translator:av_address -> CH0_YN1_L:address
	wire          ch0_yn1_l_s1_translator_avalon_anti_slave_0_chipselect;                                           // CH0_YN1_L_s1_translator:av_chipselect -> CH0_YN1_L:chipselect
	wire          ch0_yn1_l_s1_translator_avalon_anti_slave_0_write;                                                // CH0_YN1_L_s1_translator:av_write -> CH0_YN1_L:write_n
	wire   [31:0] ch0_yn1_l_s1_translator_avalon_anti_slave_0_readdata;                                             // CH0_YN1_L:readdata -> CH0_YN1_L_s1_translator:av_readdata
	wire   [31:0] ch0_yn1_ml_s1_translator_avalon_anti_slave_0_writedata;                                           // CH0_YN1_ML_s1_translator:av_writedata -> CH0_YN1_ML:writedata
	wire    [1:0] ch0_yn1_ml_s1_translator_avalon_anti_slave_0_address;                                             // CH0_YN1_ML_s1_translator:av_address -> CH0_YN1_ML:address
	wire          ch0_yn1_ml_s1_translator_avalon_anti_slave_0_chipselect;                                          // CH0_YN1_ML_s1_translator:av_chipselect -> CH0_YN1_ML:chipselect
	wire          ch0_yn1_ml_s1_translator_avalon_anti_slave_0_write;                                               // CH0_YN1_ML_s1_translator:av_write -> CH0_YN1_ML:write_n
	wire   [31:0] ch0_yn1_ml_s1_translator_avalon_anti_slave_0_readdata;                                            // CH0_YN1_ML:readdata -> CH0_YN1_ML_s1_translator:av_readdata
	wire   [31:0] ch0_yn1_mu_s1_translator_avalon_anti_slave_0_writedata;                                           // CH0_YN1_MU_s1_translator:av_writedata -> CH0_YN1_MU:writedata
	wire    [1:0] ch0_yn1_mu_s1_translator_avalon_anti_slave_0_address;                                             // CH0_YN1_MU_s1_translator:av_address -> CH0_YN1_MU:address
	wire          ch0_yn1_mu_s1_translator_avalon_anti_slave_0_chipselect;                                          // CH0_YN1_MU_s1_translator:av_chipselect -> CH0_YN1_MU:chipselect
	wire          ch0_yn1_mu_s1_translator_avalon_anti_slave_0_write;                                               // CH0_YN1_MU_s1_translator:av_write -> CH0_YN1_MU:write_n
	wire   [31:0] ch0_yn1_mu_s1_translator_avalon_anti_slave_0_readdata;                                            // CH0_YN1_MU:readdata -> CH0_YN1_MU_s1_translator:av_readdata
	wire   [31:0] ch0_yn1_u_s1_translator_avalon_anti_slave_0_writedata;                                            // CH0_YN1_U_s1_translator:av_writedata -> CH0_YN1_U:writedata
	wire    [1:0] ch0_yn1_u_s1_translator_avalon_anti_slave_0_address;                                              // CH0_YN1_U_s1_translator:av_address -> CH0_YN1_U:address
	wire          ch0_yn1_u_s1_translator_avalon_anti_slave_0_chipselect;                                           // CH0_YN1_U_s1_translator:av_chipselect -> CH0_YN1_U:chipselect
	wire          ch0_yn1_u_s1_translator_avalon_anti_slave_0_write;                                                // CH0_YN1_U_s1_translator:av_write -> CH0_YN1_U:write_n
	wire   [31:0] ch0_yn1_u_s1_translator_avalon_anti_slave_0_readdata;                                             // CH0_YN1_U:readdata -> CH0_YN1_U_s1_translator:av_readdata
	wire   [31:0] ch0_time_s1_translator_avalon_anti_slave_0_writedata;                                             // CH0_TIME_s1_translator:av_writedata -> CH0_TIME:writedata
	wire    [1:0] ch0_time_s1_translator_avalon_anti_slave_0_address;                                               // CH0_TIME_s1_translator:av_address -> CH0_TIME:address
	wire          ch0_time_s1_translator_avalon_anti_slave_0_chipselect;                                            // CH0_TIME_s1_translator:av_chipselect -> CH0_TIME:chipselect
	wire          ch0_time_s1_translator_avalon_anti_slave_0_write;                                                 // CH0_TIME_s1_translator:av_write -> CH0_TIME:write_n
	wire   [31:0] ch0_time_s1_translator_avalon_anti_slave_0_readdata;                                              // CH0_TIME:readdata -> CH0_TIME_s1_translator:av_readdata
	wire   [31:0] ch0_yn2_mu_s1_translator_avalon_anti_slave_0_writedata;                                           // CH0_YN2_MU_s1_translator:av_writedata -> CH0_YN2_MU:writedata
	wire    [1:0] ch0_yn2_mu_s1_translator_avalon_anti_slave_0_address;                                             // CH0_YN2_MU_s1_translator:av_address -> CH0_YN2_MU:address
	wire          ch0_yn2_mu_s1_translator_avalon_anti_slave_0_chipselect;                                          // CH0_YN2_MU_s1_translator:av_chipselect -> CH0_YN2_MU:chipselect
	wire          ch0_yn2_mu_s1_translator_avalon_anti_slave_0_write;                                               // CH0_YN2_MU_s1_translator:av_write -> CH0_YN2_MU:write_n
	wire   [31:0] ch0_yn2_mu_s1_translator_avalon_anti_slave_0_readdata;                                            // CH0_YN2_MU:readdata -> CH0_YN2_MU_s1_translator:av_readdata
	wire   [31:0] ch0_yn2_ml_s1_translator_avalon_anti_slave_0_writedata;                                           // CH0_YN2_ML_s1_translator:av_writedata -> CH0_YN2_ML:writedata
	wire    [1:0] ch0_yn2_ml_s1_translator_avalon_anti_slave_0_address;                                             // CH0_YN2_ML_s1_translator:av_address -> CH0_YN2_ML:address
	wire          ch0_yn2_ml_s1_translator_avalon_anti_slave_0_chipselect;                                          // CH0_YN2_ML_s1_translator:av_chipselect -> CH0_YN2_ML:chipselect
	wire          ch0_yn2_ml_s1_translator_avalon_anti_slave_0_write;                                               // CH0_YN2_ML_s1_translator:av_write -> CH0_YN2_ML:write_n
	wire   [31:0] ch0_yn2_ml_s1_translator_avalon_anti_slave_0_readdata;                                            // CH0_YN2_ML:readdata -> CH0_YN2_ML_s1_translator:av_readdata
	wire   [31:0] ch0_yn2_u_s1_translator_avalon_anti_slave_0_writedata;                                            // CH0_YN2_U_s1_translator:av_writedata -> CH0_YN2_U:writedata
	wire    [1:0] ch0_yn2_u_s1_translator_avalon_anti_slave_0_address;                                              // CH0_YN2_U_s1_translator:av_address -> CH0_YN2_U:address
	wire          ch0_yn2_u_s1_translator_avalon_anti_slave_0_chipselect;                                           // CH0_YN2_U_s1_translator:av_chipselect -> CH0_YN2_U:chipselect
	wire          ch0_yn2_u_s1_translator_avalon_anti_slave_0_write;                                                // CH0_YN2_U_s1_translator:av_write -> CH0_YN2_U:write_n
	wire   [31:0] ch0_yn2_u_s1_translator_avalon_anti_slave_0_readdata;                                             // CH0_YN2_U:readdata -> CH0_YN2_U_s1_translator:av_readdata
	wire   [31:0] ch0_yn2_l_s1_translator_avalon_anti_slave_0_writedata;                                            // CH0_YN2_L_s1_translator:av_writedata -> CH0_YN2_L:writedata
	wire    [1:0] ch0_yn2_l_s1_translator_avalon_anti_slave_0_address;                                              // CH0_YN2_L_s1_translator:av_address -> CH0_YN2_L:address
	wire          ch0_yn2_l_s1_translator_avalon_anti_slave_0_chipselect;                                           // CH0_YN2_L_s1_translator:av_chipselect -> CH0_YN2_L:chipselect
	wire          ch0_yn2_l_s1_translator_avalon_anti_slave_0_write;                                                // CH0_YN2_L_s1_translator:av_write -> CH0_YN2_L:write_n
	wire   [31:0] ch0_yn2_l_s1_translator_avalon_anti_slave_0_readdata;                                             // CH0_YN2_L:readdata -> CH0_YN2_L_s1_translator:av_readdata
	wire   [31:0] ch0_yn3_l_s1_translator_avalon_anti_slave_0_writedata;                                            // CH0_YN3_L_s1_translator:av_writedata -> CH0_YN3_L:writedata
	wire    [1:0] ch0_yn3_l_s1_translator_avalon_anti_slave_0_address;                                              // CH0_YN3_L_s1_translator:av_address -> CH0_YN3_L:address
	wire          ch0_yn3_l_s1_translator_avalon_anti_slave_0_chipselect;                                           // CH0_YN3_L_s1_translator:av_chipselect -> CH0_YN3_L:chipselect
	wire          ch0_yn3_l_s1_translator_avalon_anti_slave_0_write;                                                // CH0_YN3_L_s1_translator:av_write -> CH0_YN3_L:write_n
	wire   [31:0] ch0_yn3_l_s1_translator_avalon_anti_slave_0_readdata;                                             // CH0_YN3_L:readdata -> CH0_YN3_L_s1_translator:av_readdata
	wire   [31:0] ch0_yn3_ml_s1_translator_avalon_anti_slave_0_writedata;                                           // CH0_YN3_ML_s1_translator:av_writedata -> CH0_YN3_ML:writedata
	wire    [1:0] ch0_yn3_ml_s1_translator_avalon_anti_slave_0_address;                                             // CH0_YN3_ML_s1_translator:av_address -> CH0_YN3_ML:address
	wire          ch0_yn3_ml_s1_translator_avalon_anti_slave_0_chipselect;                                          // CH0_YN3_ML_s1_translator:av_chipselect -> CH0_YN3_ML:chipselect
	wire          ch0_yn3_ml_s1_translator_avalon_anti_slave_0_write;                                               // CH0_YN3_ML_s1_translator:av_write -> CH0_YN3_ML:write_n
	wire   [31:0] ch0_yn3_ml_s1_translator_avalon_anti_slave_0_readdata;                                            // CH0_YN3_ML:readdata -> CH0_YN3_ML_s1_translator:av_readdata
	wire   [31:0] ch0_yn3_mu_s1_translator_avalon_anti_slave_0_writedata;                                           // CH0_YN3_MU_s1_translator:av_writedata -> CH0_YN3_MU:writedata
	wire    [1:0] ch0_yn3_mu_s1_translator_avalon_anti_slave_0_address;                                             // CH0_YN3_MU_s1_translator:av_address -> CH0_YN3_MU:address
	wire          ch0_yn3_mu_s1_translator_avalon_anti_slave_0_chipselect;                                          // CH0_YN3_MU_s1_translator:av_chipselect -> CH0_YN3_MU:chipselect
	wire          ch0_yn3_mu_s1_translator_avalon_anti_slave_0_write;                                               // CH0_YN3_MU_s1_translator:av_write -> CH0_YN3_MU:write_n
	wire   [31:0] ch0_yn3_mu_s1_translator_avalon_anti_slave_0_readdata;                                            // CH0_YN3_MU:readdata -> CH0_YN3_MU_s1_translator:av_readdata
	wire   [31:0] ch0_yn3_u_s1_translator_avalon_anti_slave_0_writedata;                                            // CH0_YN3_U_s1_translator:av_writedata -> CH0_YN3_U:writedata
	wire    [1:0] ch0_yn3_u_s1_translator_avalon_anti_slave_0_address;                                              // CH0_YN3_U_s1_translator:av_address -> CH0_YN3_U:address
	wire          ch0_yn3_u_s1_translator_avalon_anti_slave_0_chipselect;                                           // CH0_YN3_U_s1_translator:av_chipselect -> CH0_YN3_U:chipselect
	wire          ch0_yn3_u_s1_translator_avalon_anti_slave_0_write;                                                // CH0_YN3_U_s1_translator:av_write -> CH0_YN3_U:write_n
	wire   [31:0] ch0_yn3_u_s1_translator_avalon_anti_slave_0_readdata;                                             // CH0_YN3_U:readdata -> CH0_YN3_U_s1_translator:av_readdata
	wire   [31:0] ch1_timer_rst_s1_translator_avalon_anti_slave_0_writedata;                                        // CH1_TIMER_RST_s1_translator:av_writedata -> CH1_TIMER_RST:writedata
	wire    [1:0] ch1_timer_rst_s1_translator_avalon_anti_slave_0_address;                                          // CH1_TIMER_RST_s1_translator:av_address -> CH1_TIMER_RST:address
	wire          ch1_timer_rst_s1_translator_avalon_anti_slave_0_chipselect;                                       // CH1_TIMER_RST_s1_translator:av_chipselect -> CH1_TIMER_RST:chipselect
	wire          ch1_timer_rst_s1_translator_avalon_anti_slave_0_write;                                            // CH1_TIMER_RST_s1_translator:av_write -> CH1_TIMER_RST:write_n
	wire   [31:0] ch1_timer_rst_s1_translator_avalon_anti_slave_0_readdata;                                         // CH1_TIMER_RST:readdata -> CH1_TIMER_RST_s1_translator:av_readdata
	wire   [31:0] ch1_thresh_s1_translator_avalon_anti_slave_0_writedata;                                           // CH1_THRESH_s1_translator:av_writedata -> CH1_THRESH:writedata
	wire    [1:0] ch1_thresh_s1_translator_avalon_anti_slave_0_address;                                             // CH1_THRESH_s1_translator:av_address -> CH1_THRESH:address
	wire          ch1_thresh_s1_translator_avalon_anti_slave_0_chipselect;                                          // CH1_THRESH_s1_translator:av_chipselect -> CH1_THRESH:chipselect
	wire          ch1_thresh_s1_translator_avalon_anti_slave_0_write;                                               // CH1_THRESH_s1_translator:av_write -> CH1_THRESH:write_n
	wire   [31:0] ch1_thresh_s1_translator_avalon_anti_slave_0_readdata;                                            // CH1_THRESH:readdata -> CH1_THRESH_s1_translator:av_readdata
	wire   [31:0] ch1_rd_peak_s1_translator_avalon_anti_slave_0_writedata;                                          // CH1_RD_PEAK_s1_translator:av_writedata -> CH1_RD_PEAK:writedata
	wire    [1:0] ch1_rd_peak_s1_translator_avalon_anti_slave_0_address;                                            // CH1_RD_PEAK_s1_translator:av_address -> CH1_RD_PEAK:address
	wire          ch1_rd_peak_s1_translator_avalon_anti_slave_0_chipselect;                                         // CH1_RD_PEAK_s1_translator:av_chipselect -> CH1_RD_PEAK:chipselect
	wire          ch1_rd_peak_s1_translator_avalon_anti_slave_0_write;                                              // CH1_RD_PEAK_s1_translator:av_write -> CH1_RD_PEAK:write_n
	wire   [31:0] ch1_rd_peak_s1_translator_avalon_anti_slave_0_readdata;                                           // CH1_RD_PEAK:readdata -> CH1_RD_PEAK_s1_translator:av_readdata
	wire   [31:0] ch1_peak_found_s1_translator_avalon_anti_slave_0_writedata;                                       // CH1_PEAK_FOUND_s1_translator:av_writedata -> CH1_PEAK_FOUND:writedata
	wire    [1:0] ch1_peak_found_s1_translator_avalon_anti_slave_0_address;                                         // CH1_PEAK_FOUND_s1_translator:av_address -> CH1_PEAK_FOUND:address
	wire          ch1_peak_found_s1_translator_avalon_anti_slave_0_chipselect;                                      // CH1_PEAK_FOUND_s1_translator:av_chipselect -> CH1_PEAK_FOUND:chipselect
	wire          ch1_peak_found_s1_translator_avalon_anti_slave_0_write;                                           // CH1_PEAK_FOUND_s1_translator:av_write -> CH1_PEAK_FOUND:write_n
	wire   [31:0] ch1_peak_found_s1_translator_avalon_anti_slave_0_readdata;                                        // CH1_PEAK_FOUND:readdata -> CH1_PEAK_FOUND_s1_translator:av_readdata
	wire   [31:0] ch1_time_s1_translator_avalon_anti_slave_0_writedata;                                             // CH1_TIME_s1_translator:av_writedata -> CH1_TIME:writedata
	wire    [1:0] ch1_time_s1_translator_avalon_anti_slave_0_address;                                               // CH1_TIME_s1_translator:av_address -> CH1_TIME:address
	wire          ch1_time_s1_translator_avalon_anti_slave_0_chipselect;                                            // CH1_TIME_s1_translator:av_chipselect -> CH1_TIME:chipselect
	wire          ch1_time_s1_translator_avalon_anti_slave_0_write;                                                 // CH1_TIME_s1_translator:av_write -> CH1_TIME:write_n
	wire   [31:0] ch1_time_s1_translator_avalon_anti_slave_0_readdata;                                              // CH1_TIME:readdata -> CH1_TIME_s1_translator:av_readdata
	wire   [31:0] ch1_yn1_u_s1_translator_avalon_anti_slave_0_writedata;                                            // CH1_YN1_U_s1_translator:av_writedata -> CH1_YN1_U:writedata
	wire    [1:0] ch1_yn1_u_s1_translator_avalon_anti_slave_0_address;                                              // CH1_YN1_U_s1_translator:av_address -> CH1_YN1_U:address
	wire          ch1_yn1_u_s1_translator_avalon_anti_slave_0_chipselect;                                           // CH1_YN1_U_s1_translator:av_chipselect -> CH1_YN1_U:chipselect
	wire          ch1_yn1_u_s1_translator_avalon_anti_slave_0_write;                                                // CH1_YN1_U_s1_translator:av_write -> CH1_YN1_U:write_n
	wire   [31:0] ch1_yn1_u_s1_translator_avalon_anti_slave_0_readdata;                                             // CH1_YN1_U:readdata -> CH1_YN1_U_s1_translator:av_readdata
	wire   [31:0] ch1_yn1_mu_s1_translator_avalon_anti_slave_0_writedata;                                           // CH1_YN1_MU_s1_translator:av_writedata -> CH1_YN1_MU:writedata
	wire    [1:0] ch1_yn1_mu_s1_translator_avalon_anti_slave_0_address;                                             // CH1_YN1_MU_s1_translator:av_address -> CH1_YN1_MU:address
	wire          ch1_yn1_mu_s1_translator_avalon_anti_slave_0_chipselect;                                          // CH1_YN1_MU_s1_translator:av_chipselect -> CH1_YN1_MU:chipselect
	wire          ch1_yn1_mu_s1_translator_avalon_anti_slave_0_write;                                               // CH1_YN1_MU_s1_translator:av_write -> CH1_YN1_MU:write_n
	wire   [31:0] ch1_yn1_mu_s1_translator_avalon_anti_slave_0_readdata;                                            // CH1_YN1_MU:readdata -> CH1_YN1_MU_s1_translator:av_readdata
	wire   [31:0] ch1_yn1_ml_s1_translator_avalon_anti_slave_0_writedata;                                           // CH1_YN1_ML_s1_translator:av_writedata -> CH1_YN1_ML:writedata
	wire    [1:0] ch1_yn1_ml_s1_translator_avalon_anti_slave_0_address;                                             // CH1_YN1_ML_s1_translator:av_address -> CH1_YN1_ML:address
	wire          ch1_yn1_ml_s1_translator_avalon_anti_slave_0_chipselect;                                          // CH1_YN1_ML_s1_translator:av_chipselect -> CH1_YN1_ML:chipselect
	wire          ch1_yn1_ml_s1_translator_avalon_anti_slave_0_write;                                               // CH1_YN1_ML_s1_translator:av_write -> CH1_YN1_ML:write_n
	wire   [31:0] ch1_yn1_ml_s1_translator_avalon_anti_slave_0_readdata;                                            // CH1_YN1_ML:readdata -> CH1_YN1_ML_s1_translator:av_readdata
	wire   [31:0] ch1_yn1_l_s1_translator_avalon_anti_slave_0_writedata;                                            // CH1_YN1_L_s1_translator:av_writedata -> CH1_YN1_L:writedata
	wire    [1:0] ch1_yn1_l_s1_translator_avalon_anti_slave_0_address;                                              // CH1_YN1_L_s1_translator:av_address -> CH1_YN1_L:address
	wire          ch1_yn1_l_s1_translator_avalon_anti_slave_0_chipselect;                                           // CH1_YN1_L_s1_translator:av_chipselect -> CH1_YN1_L:chipselect
	wire          ch1_yn1_l_s1_translator_avalon_anti_slave_0_write;                                                // CH1_YN1_L_s1_translator:av_write -> CH1_YN1_L:write_n
	wire   [31:0] ch1_yn1_l_s1_translator_avalon_anti_slave_0_readdata;                                             // CH1_YN1_L:readdata -> CH1_YN1_L_s1_translator:av_readdata
	wire   [31:0] ch1_yn2_u_s1_translator_avalon_anti_slave_0_writedata;                                            // CH1_YN2_U_s1_translator:av_writedata -> CH1_YN2_U:writedata
	wire    [1:0] ch1_yn2_u_s1_translator_avalon_anti_slave_0_address;                                              // CH1_YN2_U_s1_translator:av_address -> CH1_YN2_U:address
	wire          ch1_yn2_u_s1_translator_avalon_anti_slave_0_chipselect;                                           // CH1_YN2_U_s1_translator:av_chipselect -> CH1_YN2_U:chipselect
	wire          ch1_yn2_u_s1_translator_avalon_anti_slave_0_write;                                                // CH1_YN2_U_s1_translator:av_write -> CH1_YN2_U:write_n
	wire   [31:0] ch1_yn2_u_s1_translator_avalon_anti_slave_0_readdata;                                             // CH1_YN2_U:readdata -> CH1_YN2_U_s1_translator:av_readdata
	wire   [31:0] ch1_yn2_mu_s1_translator_avalon_anti_slave_0_writedata;                                           // CH1_YN2_MU_s1_translator:av_writedata -> CH1_YN2_MU:writedata
	wire    [1:0] ch1_yn2_mu_s1_translator_avalon_anti_slave_0_address;                                             // CH1_YN2_MU_s1_translator:av_address -> CH1_YN2_MU:address
	wire          ch1_yn2_mu_s1_translator_avalon_anti_slave_0_chipselect;                                          // CH1_YN2_MU_s1_translator:av_chipselect -> CH1_YN2_MU:chipselect
	wire          ch1_yn2_mu_s1_translator_avalon_anti_slave_0_write;                                               // CH1_YN2_MU_s1_translator:av_write -> CH1_YN2_MU:write_n
	wire   [31:0] ch1_yn2_mu_s1_translator_avalon_anti_slave_0_readdata;                                            // CH1_YN2_MU:readdata -> CH1_YN2_MU_s1_translator:av_readdata
	wire   [31:0] ch1_yn2_ml_s1_translator_avalon_anti_slave_0_writedata;                                           // CH1_YN2_ML_s1_translator:av_writedata -> CH1_YN2_ML:writedata
	wire    [1:0] ch1_yn2_ml_s1_translator_avalon_anti_slave_0_address;                                             // CH1_YN2_ML_s1_translator:av_address -> CH1_YN2_ML:address
	wire          ch1_yn2_ml_s1_translator_avalon_anti_slave_0_chipselect;                                          // CH1_YN2_ML_s1_translator:av_chipselect -> CH1_YN2_ML:chipselect
	wire          ch1_yn2_ml_s1_translator_avalon_anti_slave_0_write;                                               // CH1_YN2_ML_s1_translator:av_write -> CH1_YN2_ML:write_n
	wire   [31:0] ch1_yn2_ml_s1_translator_avalon_anti_slave_0_readdata;                                            // CH1_YN2_ML:readdata -> CH1_YN2_ML_s1_translator:av_readdata
	wire   [31:0] ch1_yn2_l_s1_translator_avalon_anti_slave_0_writedata;                                            // CH1_YN2_L_s1_translator:av_writedata -> CH1_YN2_L:writedata
	wire    [1:0] ch1_yn2_l_s1_translator_avalon_anti_slave_0_address;                                              // CH1_YN2_L_s1_translator:av_address -> CH1_YN2_L:address
	wire          ch1_yn2_l_s1_translator_avalon_anti_slave_0_chipselect;                                           // CH1_YN2_L_s1_translator:av_chipselect -> CH1_YN2_L:chipselect
	wire          ch1_yn2_l_s1_translator_avalon_anti_slave_0_write;                                                // CH1_YN2_L_s1_translator:av_write -> CH1_YN2_L:write_n
	wire   [31:0] ch1_yn2_l_s1_translator_avalon_anti_slave_0_readdata;                                             // CH1_YN2_L:readdata -> CH1_YN2_L_s1_translator:av_readdata
	wire   [31:0] ch1_yn3_u_s1_translator_avalon_anti_slave_0_writedata;                                            // CH1_YN3_U_s1_translator:av_writedata -> CH1_YN3_U:writedata
	wire    [1:0] ch1_yn3_u_s1_translator_avalon_anti_slave_0_address;                                              // CH1_YN3_U_s1_translator:av_address -> CH1_YN3_U:address
	wire          ch1_yn3_u_s1_translator_avalon_anti_slave_0_chipselect;                                           // CH1_YN3_U_s1_translator:av_chipselect -> CH1_YN3_U:chipselect
	wire          ch1_yn3_u_s1_translator_avalon_anti_slave_0_write;                                                // CH1_YN3_U_s1_translator:av_write -> CH1_YN3_U:write_n
	wire   [31:0] ch1_yn3_u_s1_translator_avalon_anti_slave_0_readdata;                                             // CH1_YN3_U:readdata -> CH1_YN3_U_s1_translator:av_readdata
	wire   [31:0] ch1_yn3_mu_s1_translator_avalon_anti_slave_0_writedata;                                           // CH1_YN3_MU_s1_translator:av_writedata -> CH1_YN3_MU:writedata
	wire    [1:0] ch1_yn3_mu_s1_translator_avalon_anti_slave_0_address;                                             // CH1_YN3_MU_s1_translator:av_address -> CH1_YN3_MU:address
	wire          ch1_yn3_mu_s1_translator_avalon_anti_slave_0_chipselect;                                          // CH1_YN3_MU_s1_translator:av_chipselect -> CH1_YN3_MU:chipselect
	wire          ch1_yn3_mu_s1_translator_avalon_anti_slave_0_write;                                               // CH1_YN3_MU_s1_translator:av_write -> CH1_YN3_MU:write_n
	wire   [31:0] ch1_yn3_mu_s1_translator_avalon_anti_slave_0_readdata;                                            // CH1_YN3_MU:readdata -> CH1_YN3_MU_s1_translator:av_readdata
	wire   [31:0] ch1_yn3_ml_s1_translator_avalon_anti_slave_0_writedata;                                           // CH1_YN3_ML_s1_translator:av_writedata -> CH1_YN3_ML:writedata
	wire    [1:0] ch1_yn3_ml_s1_translator_avalon_anti_slave_0_address;                                             // CH1_YN3_ML_s1_translator:av_address -> CH1_YN3_ML:address
	wire          ch1_yn3_ml_s1_translator_avalon_anti_slave_0_chipselect;                                          // CH1_YN3_ML_s1_translator:av_chipselect -> CH1_YN3_ML:chipselect
	wire          ch1_yn3_ml_s1_translator_avalon_anti_slave_0_write;                                               // CH1_YN3_ML_s1_translator:av_write -> CH1_YN3_ML:write_n
	wire   [31:0] ch1_yn3_ml_s1_translator_avalon_anti_slave_0_readdata;                                            // CH1_YN3_ML:readdata -> CH1_YN3_ML_s1_translator:av_readdata
	wire   [31:0] ch1_yn3_l_s1_translator_avalon_anti_slave_0_writedata;                                            // CH1_YN3_L_s1_translator:av_writedata -> CH1_YN3_L:writedata
	wire    [1:0] ch1_yn3_l_s1_translator_avalon_anti_slave_0_address;                                              // CH1_YN3_L_s1_translator:av_address -> CH1_YN3_L:address
	wire          ch1_yn3_l_s1_translator_avalon_anti_slave_0_chipselect;                                           // CH1_YN3_L_s1_translator:av_chipselect -> CH1_YN3_L:chipselect
	wire          ch1_yn3_l_s1_translator_avalon_anti_slave_0_write;                                                // CH1_YN3_L_s1_translator:av_write -> CH1_YN3_L:write_n
	wire   [31:0] ch1_yn3_l_s1_translator_avalon_anti_slave_0_readdata;                                             // CH1_YN3_L:readdata -> CH1_YN3_L_s1_translator:av_readdata
	wire   [31:0] ch2_timer_rst_s1_translator_avalon_anti_slave_0_writedata;                                        // CH2_TIMER_RST_s1_translator:av_writedata -> CH2_TIMER_RST:writedata
	wire    [1:0] ch2_timer_rst_s1_translator_avalon_anti_slave_0_address;                                          // CH2_TIMER_RST_s1_translator:av_address -> CH2_TIMER_RST:address
	wire          ch2_timer_rst_s1_translator_avalon_anti_slave_0_chipselect;                                       // CH2_TIMER_RST_s1_translator:av_chipselect -> CH2_TIMER_RST:chipselect
	wire          ch2_timer_rst_s1_translator_avalon_anti_slave_0_write;                                            // CH2_TIMER_RST_s1_translator:av_write -> CH2_TIMER_RST:write_n
	wire   [31:0] ch2_timer_rst_s1_translator_avalon_anti_slave_0_readdata;                                         // CH2_TIMER_RST:readdata -> CH2_TIMER_RST_s1_translator:av_readdata
	wire   [31:0] ch2_thresh_s1_translator_avalon_anti_slave_0_writedata;                                           // CH2_THRESH_s1_translator:av_writedata -> CH2_THRESH:writedata
	wire    [1:0] ch2_thresh_s1_translator_avalon_anti_slave_0_address;                                             // CH2_THRESH_s1_translator:av_address -> CH2_THRESH:address
	wire          ch2_thresh_s1_translator_avalon_anti_slave_0_chipselect;                                          // CH2_THRESH_s1_translator:av_chipselect -> CH2_THRESH:chipselect
	wire          ch2_thresh_s1_translator_avalon_anti_slave_0_write;                                               // CH2_THRESH_s1_translator:av_write -> CH2_THRESH:write_n
	wire   [31:0] ch2_thresh_s1_translator_avalon_anti_slave_0_readdata;                                            // CH2_THRESH:readdata -> CH2_THRESH_s1_translator:av_readdata
	wire   [31:0] ch2_rd_peak_s1_translator_avalon_anti_slave_0_writedata;                                          // CH2_RD_PEAK_s1_translator:av_writedata -> CH2_RD_PEAK:writedata
	wire    [1:0] ch2_rd_peak_s1_translator_avalon_anti_slave_0_address;                                            // CH2_RD_PEAK_s1_translator:av_address -> CH2_RD_PEAK:address
	wire          ch2_rd_peak_s1_translator_avalon_anti_slave_0_chipselect;                                         // CH2_RD_PEAK_s1_translator:av_chipselect -> CH2_RD_PEAK:chipselect
	wire          ch2_rd_peak_s1_translator_avalon_anti_slave_0_write;                                              // CH2_RD_PEAK_s1_translator:av_write -> CH2_RD_PEAK:write_n
	wire   [31:0] ch2_rd_peak_s1_translator_avalon_anti_slave_0_readdata;                                           // CH2_RD_PEAK:readdata -> CH2_RD_PEAK_s1_translator:av_readdata
	wire   [31:0] ch2_peak_found_s1_translator_avalon_anti_slave_0_writedata;                                       // CH2_PEAK_FOUND_s1_translator:av_writedata -> CH2_PEAK_FOUND:writedata
	wire    [1:0] ch2_peak_found_s1_translator_avalon_anti_slave_0_address;                                         // CH2_PEAK_FOUND_s1_translator:av_address -> CH2_PEAK_FOUND:address
	wire          ch2_peak_found_s1_translator_avalon_anti_slave_0_chipselect;                                      // CH2_PEAK_FOUND_s1_translator:av_chipselect -> CH2_PEAK_FOUND:chipselect
	wire          ch2_peak_found_s1_translator_avalon_anti_slave_0_write;                                           // CH2_PEAK_FOUND_s1_translator:av_write -> CH2_PEAK_FOUND:write_n
	wire   [31:0] ch2_peak_found_s1_translator_avalon_anti_slave_0_readdata;                                        // CH2_PEAK_FOUND:readdata -> CH2_PEAK_FOUND_s1_translator:av_readdata
	wire   [31:0] ch2_time_s1_translator_avalon_anti_slave_0_writedata;                                             // CH2_TIME_s1_translator:av_writedata -> CH2_TIME:writedata
	wire    [1:0] ch2_time_s1_translator_avalon_anti_slave_0_address;                                               // CH2_TIME_s1_translator:av_address -> CH2_TIME:address
	wire          ch2_time_s1_translator_avalon_anti_slave_0_chipselect;                                            // CH2_TIME_s1_translator:av_chipselect -> CH2_TIME:chipselect
	wire          ch2_time_s1_translator_avalon_anti_slave_0_write;                                                 // CH2_TIME_s1_translator:av_write -> CH2_TIME:write_n
	wire   [31:0] ch2_time_s1_translator_avalon_anti_slave_0_readdata;                                              // CH2_TIME:readdata -> CH2_TIME_s1_translator:av_readdata
	wire   [31:0] ch2_yn1_u_s1_translator_avalon_anti_slave_0_writedata;                                            // CH2_YN1_U_s1_translator:av_writedata -> CH2_YN1_U:writedata
	wire    [1:0] ch2_yn1_u_s1_translator_avalon_anti_slave_0_address;                                              // CH2_YN1_U_s1_translator:av_address -> CH2_YN1_U:address
	wire          ch2_yn1_u_s1_translator_avalon_anti_slave_0_chipselect;                                           // CH2_YN1_U_s1_translator:av_chipselect -> CH2_YN1_U:chipselect
	wire          ch2_yn1_u_s1_translator_avalon_anti_slave_0_write;                                                // CH2_YN1_U_s1_translator:av_write -> CH2_YN1_U:write_n
	wire   [31:0] ch2_yn1_u_s1_translator_avalon_anti_slave_0_readdata;                                             // CH2_YN1_U:readdata -> CH2_YN1_U_s1_translator:av_readdata
	wire   [31:0] ch2_yn1_mu_s1_translator_avalon_anti_slave_0_writedata;                                           // CH2_YN1_MU_s1_translator:av_writedata -> CH2_YN1_MU:writedata
	wire    [1:0] ch2_yn1_mu_s1_translator_avalon_anti_slave_0_address;                                             // CH2_YN1_MU_s1_translator:av_address -> CH2_YN1_MU:address
	wire          ch2_yn1_mu_s1_translator_avalon_anti_slave_0_chipselect;                                          // CH2_YN1_MU_s1_translator:av_chipselect -> CH2_YN1_MU:chipselect
	wire          ch2_yn1_mu_s1_translator_avalon_anti_slave_0_write;                                               // CH2_YN1_MU_s1_translator:av_write -> CH2_YN1_MU:write_n
	wire   [31:0] ch2_yn1_mu_s1_translator_avalon_anti_slave_0_readdata;                                            // CH2_YN1_MU:readdata -> CH2_YN1_MU_s1_translator:av_readdata
	wire   [31:0] ch2_yn1_ml_s1_translator_avalon_anti_slave_0_writedata;                                           // CH2_YN1_ML_s1_translator:av_writedata -> CH2_YN1_ML:writedata
	wire    [1:0] ch2_yn1_ml_s1_translator_avalon_anti_slave_0_address;                                             // CH2_YN1_ML_s1_translator:av_address -> CH2_YN1_ML:address
	wire          ch2_yn1_ml_s1_translator_avalon_anti_slave_0_chipselect;                                          // CH2_YN1_ML_s1_translator:av_chipselect -> CH2_YN1_ML:chipselect
	wire          ch2_yn1_ml_s1_translator_avalon_anti_slave_0_write;                                               // CH2_YN1_ML_s1_translator:av_write -> CH2_YN1_ML:write_n
	wire   [31:0] ch2_yn1_ml_s1_translator_avalon_anti_slave_0_readdata;                                            // CH2_YN1_ML:readdata -> CH2_YN1_ML_s1_translator:av_readdata
	wire   [31:0] ch2_yn1_l_s1_translator_avalon_anti_slave_0_writedata;                                            // CH2_YN1_L_s1_translator:av_writedata -> CH2_YN1_L:writedata
	wire    [1:0] ch2_yn1_l_s1_translator_avalon_anti_slave_0_address;                                              // CH2_YN1_L_s1_translator:av_address -> CH2_YN1_L:address
	wire          ch2_yn1_l_s1_translator_avalon_anti_slave_0_chipselect;                                           // CH2_YN1_L_s1_translator:av_chipselect -> CH2_YN1_L:chipselect
	wire          ch2_yn1_l_s1_translator_avalon_anti_slave_0_write;                                                // CH2_YN1_L_s1_translator:av_write -> CH2_YN1_L:write_n
	wire   [31:0] ch2_yn1_l_s1_translator_avalon_anti_slave_0_readdata;                                             // CH2_YN1_L:readdata -> CH2_YN1_L_s1_translator:av_readdata
	wire   [31:0] ch2_yn2_u_s1_translator_avalon_anti_slave_0_writedata;                                            // CH2_YN2_U_s1_translator:av_writedata -> CH2_YN2_U:writedata
	wire    [1:0] ch2_yn2_u_s1_translator_avalon_anti_slave_0_address;                                              // CH2_YN2_U_s1_translator:av_address -> CH2_YN2_U:address
	wire          ch2_yn2_u_s1_translator_avalon_anti_slave_0_chipselect;                                           // CH2_YN2_U_s1_translator:av_chipselect -> CH2_YN2_U:chipselect
	wire          ch2_yn2_u_s1_translator_avalon_anti_slave_0_write;                                                // CH2_YN2_U_s1_translator:av_write -> CH2_YN2_U:write_n
	wire   [31:0] ch2_yn2_u_s1_translator_avalon_anti_slave_0_readdata;                                             // CH2_YN2_U:readdata -> CH2_YN2_U_s1_translator:av_readdata
	wire   [31:0] ch2_yn2_mu_s1_translator_avalon_anti_slave_0_writedata;                                           // CH2_YN2_MU_s1_translator:av_writedata -> CH2_YN2_MU:writedata
	wire    [1:0] ch2_yn2_mu_s1_translator_avalon_anti_slave_0_address;                                             // CH2_YN2_MU_s1_translator:av_address -> CH2_YN2_MU:address
	wire          ch2_yn2_mu_s1_translator_avalon_anti_slave_0_chipselect;                                          // CH2_YN2_MU_s1_translator:av_chipselect -> CH2_YN2_MU:chipselect
	wire          ch2_yn2_mu_s1_translator_avalon_anti_slave_0_write;                                               // CH2_YN2_MU_s1_translator:av_write -> CH2_YN2_MU:write_n
	wire   [31:0] ch2_yn2_mu_s1_translator_avalon_anti_slave_0_readdata;                                            // CH2_YN2_MU:readdata -> CH2_YN2_MU_s1_translator:av_readdata
	wire   [31:0] ch2_yn2_ml_s1_translator_avalon_anti_slave_0_writedata;                                           // CH2_YN2_ML_s1_translator:av_writedata -> CH2_YN2_ML:writedata
	wire    [1:0] ch2_yn2_ml_s1_translator_avalon_anti_slave_0_address;                                             // CH2_YN2_ML_s1_translator:av_address -> CH2_YN2_ML:address
	wire          ch2_yn2_ml_s1_translator_avalon_anti_slave_0_chipselect;                                          // CH2_YN2_ML_s1_translator:av_chipselect -> CH2_YN2_ML:chipselect
	wire          ch2_yn2_ml_s1_translator_avalon_anti_slave_0_write;                                               // CH2_YN2_ML_s1_translator:av_write -> CH2_YN2_ML:write_n
	wire   [31:0] ch2_yn2_ml_s1_translator_avalon_anti_slave_0_readdata;                                            // CH2_YN2_ML:readdata -> CH2_YN2_ML_s1_translator:av_readdata
	wire   [31:0] ch2_yn2_l_s1_translator_avalon_anti_slave_0_writedata;                                            // CH2_YN2_L_s1_translator:av_writedata -> CH2_YN2_L:writedata
	wire    [1:0] ch2_yn2_l_s1_translator_avalon_anti_slave_0_address;                                              // CH2_YN2_L_s1_translator:av_address -> CH2_YN2_L:address
	wire          ch2_yn2_l_s1_translator_avalon_anti_slave_0_chipselect;                                           // CH2_YN2_L_s1_translator:av_chipselect -> CH2_YN2_L:chipselect
	wire          ch2_yn2_l_s1_translator_avalon_anti_slave_0_write;                                                // CH2_YN2_L_s1_translator:av_write -> CH2_YN2_L:write_n
	wire   [31:0] ch2_yn2_l_s1_translator_avalon_anti_slave_0_readdata;                                             // CH2_YN2_L:readdata -> CH2_YN2_L_s1_translator:av_readdata
	wire   [31:0] ch2_yn3_u_s1_translator_avalon_anti_slave_0_writedata;                                            // CH2_YN3_U_s1_translator:av_writedata -> CH2_YN3_U:writedata
	wire    [1:0] ch2_yn3_u_s1_translator_avalon_anti_slave_0_address;                                              // CH2_YN3_U_s1_translator:av_address -> CH2_YN3_U:address
	wire          ch2_yn3_u_s1_translator_avalon_anti_slave_0_chipselect;                                           // CH2_YN3_U_s1_translator:av_chipselect -> CH2_YN3_U:chipselect
	wire          ch2_yn3_u_s1_translator_avalon_anti_slave_0_write;                                                // CH2_YN3_U_s1_translator:av_write -> CH2_YN3_U:write_n
	wire   [31:0] ch2_yn3_u_s1_translator_avalon_anti_slave_0_readdata;                                             // CH2_YN3_U:readdata -> CH2_YN3_U_s1_translator:av_readdata
	wire   [31:0] ch2_yn3_mu_s1_translator_avalon_anti_slave_0_writedata;                                           // CH2_YN3_MU_s1_translator:av_writedata -> CH2_YN3_MU:writedata
	wire    [1:0] ch2_yn3_mu_s1_translator_avalon_anti_slave_0_address;                                             // CH2_YN3_MU_s1_translator:av_address -> CH2_YN3_MU:address
	wire          ch2_yn3_mu_s1_translator_avalon_anti_slave_0_chipselect;                                          // CH2_YN3_MU_s1_translator:av_chipselect -> CH2_YN3_MU:chipselect
	wire          ch2_yn3_mu_s1_translator_avalon_anti_slave_0_write;                                               // CH2_YN3_MU_s1_translator:av_write -> CH2_YN3_MU:write_n
	wire   [31:0] ch2_yn3_mu_s1_translator_avalon_anti_slave_0_readdata;                                            // CH2_YN3_MU:readdata -> CH2_YN3_MU_s1_translator:av_readdata
	wire   [31:0] ch2_yn3_ml_s1_translator_avalon_anti_slave_0_writedata;                                           // CH2_YN3_ML_s1_translator:av_writedata -> CH2_YN3_ML:writedata
	wire    [1:0] ch2_yn3_ml_s1_translator_avalon_anti_slave_0_address;                                             // CH2_YN3_ML_s1_translator:av_address -> CH2_YN3_ML:address
	wire          ch2_yn3_ml_s1_translator_avalon_anti_slave_0_chipselect;                                          // CH2_YN3_ML_s1_translator:av_chipselect -> CH2_YN3_ML:chipselect
	wire          ch2_yn3_ml_s1_translator_avalon_anti_slave_0_write;                                               // CH2_YN3_ML_s1_translator:av_write -> CH2_YN3_ML:write_n
	wire   [31:0] ch2_yn3_ml_s1_translator_avalon_anti_slave_0_readdata;                                            // CH2_YN3_ML:readdata -> CH2_YN3_ML_s1_translator:av_readdata
	wire   [31:0] ch2_yn3_l_s1_translator_avalon_anti_slave_0_writedata;                                            // CH2_YN3_L_s1_translator:av_writedata -> CH2_YN3_L:writedata
	wire    [1:0] ch2_yn3_l_s1_translator_avalon_anti_slave_0_address;                                              // CH2_YN3_L_s1_translator:av_address -> CH2_YN3_L:address
	wire          ch2_yn3_l_s1_translator_avalon_anti_slave_0_chipselect;                                           // CH2_YN3_L_s1_translator:av_chipselect -> CH2_YN3_L:chipselect
	wire          ch2_yn3_l_s1_translator_avalon_anti_slave_0_write;                                                // CH2_YN3_L_s1_translator:av_write -> CH2_YN3_L:write_n
	wire   [31:0] ch2_yn3_l_s1_translator_avalon_anti_slave_0_readdata;                                             // CH2_YN3_L:readdata -> CH2_YN3_L_s1_translator:av_readdata
	wire   [31:0] ch3_timer_rst_s1_translator_avalon_anti_slave_0_writedata;                                        // CH3_TIMER_RST_s1_translator:av_writedata -> CH3_TIMER_RST:writedata
	wire    [1:0] ch3_timer_rst_s1_translator_avalon_anti_slave_0_address;                                          // CH3_TIMER_RST_s1_translator:av_address -> CH3_TIMER_RST:address
	wire          ch3_timer_rst_s1_translator_avalon_anti_slave_0_chipselect;                                       // CH3_TIMER_RST_s1_translator:av_chipselect -> CH3_TIMER_RST:chipselect
	wire          ch3_timer_rst_s1_translator_avalon_anti_slave_0_write;                                            // CH3_TIMER_RST_s1_translator:av_write -> CH3_TIMER_RST:write_n
	wire   [31:0] ch3_timer_rst_s1_translator_avalon_anti_slave_0_readdata;                                         // CH3_TIMER_RST:readdata -> CH3_TIMER_RST_s1_translator:av_readdata
	wire   [31:0] ch3_thresh_s1_translator_avalon_anti_slave_0_writedata;                                           // CH3_THRESH_s1_translator:av_writedata -> CH3_THRESH:writedata
	wire    [1:0] ch3_thresh_s1_translator_avalon_anti_slave_0_address;                                             // CH3_THRESH_s1_translator:av_address -> CH3_THRESH:address
	wire          ch3_thresh_s1_translator_avalon_anti_slave_0_chipselect;                                          // CH3_THRESH_s1_translator:av_chipselect -> CH3_THRESH:chipselect
	wire          ch3_thresh_s1_translator_avalon_anti_slave_0_write;                                               // CH3_THRESH_s1_translator:av_write -> CH3_THRESH:write_n
	wire   [31:0] ch3_thresh_s1_translator_avalon_anti_slave_0_readdata;                                            // CH3_THRESH:readdata -> CH3_THRESH_s1_translator:av_readdata
	wire   [31:0] ch3_rd_peak_s1_translator_avalon_anti_slave_0_writedata;                                          // CH3_RD_PEAK_s1_translator:av_writedata -> CH3_RD_PEAK:writedata
	wire    [1:0] ch3_rd_peak_s1_translator_avalon_anti_slave_0_address;                                            // CH3_RD_PEAK_s1_translator:av_address -> CH3_RD_PEAK:address
	wire          ch3_rd_peak_s1_translator_avalon_anti_slave_0_chipselect;                                         // CH3_RD_PEAK_s1_translator:av_chipselect -> CH3_RD_PEAK:chipselect
	wire          ch3_rd_peak_s1_translator_avalon_anti_slave_0_write;                                              // CH3_RD_PEAK_s1_translator:av_write -> CH3_RD_PEAK:write_n
	wire   [31:0] ch3_rd_peak_s1_translator_avalon_anti_slave_0_readdata;                                           // CH3_RD_PEAK:readdata -> CH3_RD_PEAK_s1_translator:av_readdata
	wire   [31:0] ch3_peak_found_s1_translator_avalon_anti_slave_0_writedata;                                       // CH3_PEAK_FOUND_s1_translator:av_writedata -> CH3_PEAK_FOUND:writedata
	wire    [1:0] ch3_peak_found_s1_translator_avalon_anti_slave_0_address;                                         // CH3_PEAK_FOUND_s1_translator:av_address -> CH3_PEAK_FOUND:address
	wire          ch3_peak_found_s1_translator_avalon_anti_slave_0_chipselect;                                      // CH3_PEAK_FOUND_s1_translator:av_chipselect -> CH3_PEAK_FOUND:chipselect
	wire          ch3_peak_found_s1_translator_avalon_anti_slave_0_write;                                           // CH3_PEAK_FOUND_s1_translator:av_write -> CH3_PEAK_FOUND:write_n
	wire   [31:0] ch3_peak_found_s1_translator_avalon_anti_slave_0_readdata;                                        // CH3_PEAK_FOUND:readdata -> CH3_PEAK_FOUND_s1_translator:av_readdata
	wire   [31:0] ch3_yn1_u_s1_translator_avalon_anti_slave_0_writedata;                                            // CH3_YN1_U_s1_translator:av_writedata -> CH3_YN1_U:writedata
	wire    [1:0] ch3_yn1_u_s1_translator_avalon_anti_slave_0_address;                                              // CH3_YN1_U_s1_translator:av_address -> CH3_YN1_U:address
	wire          ch3_yn1_u_s1_translator_avalon_anti_slave_0_chipselect;                                           // CH3_YN1_U_s1_translator:av_chipselect -> CH3_YN1_U:chipselect
	wire          ch3_yn1_u_s1_translator_avalon_anti_slave_0_write;                                                // CH3_YN1_U_s1_translator:av_write -> CH3_YN1_U:write_n
	wire   [31:0] ch3_yn1_u_s1_translator_avalon_anti_slave_0_readdata;                                             // CH3_YN1_U:readdata -> CH3_YN1_U_s1_translator:av_readdata
	wire   [31:0] ch3_time_s1_translator_avalon_anti_slave_0_writedata;                                             // CH3_TIME_s1_translator:av_writedata -> CH3_TIME:writedata
	wire    [1:0] ch3_time_s1_translator_avalon_anti_slave_0_address;                                               // CH3_TIME_s1_translator:av_address -> CH3_TIME:address
	wire          ch3_time_s1_translator_avalon_anti_slave_0_chipselect;                                            // CH3_TIME_s1_translator:av_chipselect -> CH3_TIME:chipselect
	wire          ch3_time_s1_translator_avalon_anti_slave_0_write;                                                 // CH3_TIME_s1_translator:av_write -> CH3_TIME:write_n
	wire   [31:0] ch3_time_s1_translator_avalon_anti_slave_0_readdata;                                              // CH3_TIME:readdata -> CH3_TIME_s1_translator:av_readdata
	wire   [31:0] ch3_yn3_l_s1_translator_avalon_anti_slave_0_writedata;                                            // CH3_YN3_L_s1_translator:av_writedata -> CH3_YN3_L:writedata
	wire    [1:0] ch3_yn3_l_s1_translator_avalon_anti_slave_0_address;                                              // CH3_YN3_L_s1_translator:av_address -> CH3_YN3_L:address
	wire          ch3_yn3_l_s1_translator_avalon_anti_slave_0_chipselect;                                           // CH3_YN3_L_s1_translator:av_chipselect -> CH3_YN3_L:chipselect
	wire          ch3_yn3_l_s1_translator_avalon_anti_slave_0_write;                                                // CH3_YN3_L_s1_translator:av_write -> CH3_YN3_L:write_n
	wire   [31:0] ch3_yn3_l_s1_translator_avalon_anti_slave_0_readdata;                                             // CH3_YN3_L:readdata -> CH3_YN3_L_s1_translator:av_readdata
	wire   [31:0] ch3_yn3_ml_s1_translator_avalon_anti_slave_0_writedata;                                           // CH3_YN3_ML_s1_translator:av_writedata -> CH3_YN3_ML:writedata
	wire    [1:0] ch3_yn3_ml_s1_translator_avalon_anti_slave_0_address;                                             // CH3_YN3_ML_s1_translator:av_address -> CH3_YN3_ML:address
	wire          ch3_yn3_ml_s1_translator_avalon_anti_slave_0_chipselect;                                          // CH3_YN3_ML_s1_translator:av_chipselect -> CH3_YN3_ML:chipselect
	wire          ch3_yn3_ml_s1_translator_avalon_anti_slave_0_write;                                               // CH3_YN3_ML_s1_translator:av_write -> CH3_YN3_ML:write_n
	wire   [31:0] ch3_yn3_ml_s1_translator_avalon_anti_slave_0_readdata;                                            // CH3_YN3_ML:readdata -> CH3_YN3_ML_s1_translator:av_readdata
	wire   [31:0] ch3_yn3_mu_s1_translator_avalon_anti_slave_0_writedata;                                           // CH3_YN3_MU_s1_translator:av_writedata -> CH3_YN3_MU:writedata
	wire    [1:0] ch3_yn3_mu_s1_translator_avalon_anti_slave_0_address;                                             // CH3_YN3_MU_s1_translator:av_address -> CH3_YN3_MU:address
	wire          ch3_yn3_mu_s1_translator_avalon_anti_slave_0_chipselect;                                          // CH3_YN3_MU_s1_translator:av_chipselect -> CH3_YN3_MU:chipselect
	wire          ch3_yn3_mu_s1_translator_avalon_anti_slave_0_write;                                               // CH3_YN3_MU_s1_translator:av_write -> CH3_YN3_MU:write_n
	wire   [31:0] ch3_yn3_mu_s1_translator_avalon_anti_slave_0_readdata;                                            // CH3_YN3_MU:readdata -> CH3_YN3_MU_s1_translator:av_readdata
	wire   [31:0] ch3_yn3_u_s1_translator_avalon_anti_slave_0_writedata;                                            // CH3_YN3_U_s1_translator:av_writedata -> CH3_YN3_U:writedata
	wire    [1:0] ch3_yn3_u_s1_translator_avalon_anti_slave_0_address;                                              // CH3_YN3_U_s1_translator:av_address -> CH3_YN3_U:address
	wire          ch3_yn3_u_s1_translator_avalon_anti_slave_0_chipselect;                                           // CH3_YN3_U_s1_translator:av_chipselect -> CH3_YN3_U:chipselect
	wire          ch3_yn3_u_s1_translator_avalon_anti_slave_0_write;                                                // CH3_YN3_U_s1_translator:av_write -> CH3_YN3_U:write_n
	wire   [31:0] ch3_yn3_u_s1_translator_avalon_anti_slave_0_readdata;                                             // CH3_YN3_U:readdata -> CH3_YN3_U_s1_translator:av_readdata
	wire   [31:0] ch3_yn2_l_s1_translator_avalon_anti_slave_0_writedata;                                            // CH3_YN2_L_s1_translator:av_writedata -> CH3_YN2_L:writedata
	wire    [1:0] ch3_yn2_l_s1_translator_avalon_anti_slave_0_address;                                              // CH3_YN2_L_s1_translator:av_address -> CH3_YN2_L:address
	wire          ch3_yn2_l_s1_translator_avalon_anti_slave_0_chipselect;                                           // CH3_YN2_L_s1_translator:av_chipselect -> CH3_YN2_L:chipselect
	wire          ch3_yn2_l_s1_translator_avalon_anti_slave_0_write;                                                // CH3_YN2_L_s1_translator:av_write -> CH3_YN2_L:write_n
	wire   [31:0] ch3_yn2_l_s1_translator_avalon_anti_slave_0_readdata;                                             // CH3_YN2_L:readdata -> CH3_YN2_L_s1_translator:av_readdata
	wire   [31:0] ch3_yn2_ml_s1_translator_avalon_anti_slave_0_writedata;                                           // CH3_YN2_ML_s1_translator:av_writedata -> CH3_YN2_ML:writedata
	wire    [1:0] ch3_yn2_ml_s1_translator_avalon_anti_slave_0_address;                                             // CH3_YN2_ML_s1_translator:av_address -> CH3_YN2_ML:address
	wire          ch3_yn2_ml_s1_translator_avalon_anti_slave_0_chipselect;                                          // CH3_YN2_ML_s1_translator:av_chipselect -> CH3_YN2_ML:chipselect
	wire          ch3_yn2_ml_s1_translator_avalon_anti_slave_0_write;                                               // CH3_YN2_ML_s1_translator:av_write -> CH3_YN2_ML:write_n
	wire   [31:0] ch3_yn2_ml_s1_translator_avalon_anti_slave_0_readdata;                                            // CH3_YN2_ML:readdata -> CH3_YN2_ML_s1_translator:av_readdata
	wire   [31:0] ch3_yn2_mu_s1_translator_avalon_anti_slave_0_writedata;                                           // CH3_YN2_MU_s1_translator:av_writedata -> CH3_YN2_MU:writedata
	wire    [1:0] ch3_yn2_mu_s1_translator_avalon_anti_slave_0_address;                                             // CH3_YN2_MU_s1_translator:av_address -> CH3_YN2_MU:address
	wire          ch3_yn2_mu_s1_translator_avalon_anti_slave_0_chipselect;                                          // CH3_YN2_MU_s1_translator:av_chipselect -> CH3_YN2_MU:chipselect
	wire          ch3_yn2_mu_s1_translator_avalon_anti_slave_0_write;                                               // CH3_YN2_MU_s1_translator:av_write -> CH3_YN2_MU:write_n
	wire   [31:0] ch3_yn2_mu_s1_translator_avalon_anti_slave_0_readdata;                                            // CH3_YN2_MU:readdata -> CH3_YN2_MU_s1_translator:av_readdata
	wire   [31:0] ch3_yn2_u_s1_translator_avalon_anti_slave_0_writedata;                                            // CH3_YN2_U_s1_translator:av_writedata -> CH3_YN2_U:writedata
	wire    [1:0] ch3_yn2_u_s1_translator_avalon_anti_slave_0_address;                                              // CH3_YN2_U_s1_translator:av_address -> CH3_YN2_U:address
	wire          ch3_yn2_u_s1_translator_avalon_anti_slave_0_chipselect;                                           // CH3_YN2_U_s1_translator:av_chipselect -> CH3_YN2_U:chipselect
	wire          ch3_yn2_u_s1_translator_avalon_anti_slave_0_write;                                                // CH3_YN2_U_s1_translator:av_write -> CH3_YN2_U:write_n
	wire   [31:0] ch3_yn2_u_s1_translator_avalon_anti_slave_0_readdata;                                             // CH3_YN2_U:readdata -> CH3_YN2_U_s1_translator:av_readdata
	wire   [31:0] ch3_yn1_l_s1_translator_avalon_anti_slave_0_writedata;                                            // CH3_YN1_L_s1_translator:av_writedata -> CH3_YN1_L:writedata
	wire    [1:0] ch3_yn1_l_s1_translator_avalon_anti_slave_0_address;                                              // CH3_YN1_L_s1_translator:av_address -> CH3_YN1_L:address
	wire          ch3_yn1_l_s1_translator_avalon_anti_slave_0_chipselect;                                           // CH3_YN1_L_s1_translator:av_chipselect -> CH3_YN1_L:chipselect
	wire          ch3_yn1_l_s1_translator_avalon_anti_slave_0_write;                                                // CH3_YN1_L_s1_translator:av_write -> CH3_YN1_L:write_n
	wire   [31:0] ch3_yn1_l_s1_translator_avalon_anti_slave_0_readdata;                                             // CH3_YN1_L:readdata -> CH3_YN1_L_s1_translator:av_readdata
	wire   [31:0] ch3_yn1_mu_s1_translator_avalon_anti_slave_0_writedata;                                           // CH3_YN1_MU_s1_translator:av_writedata -> CH3_YN1_MU:writedata
	wire    [1:0] ch3_yn1_mu_s1_translator_avalon_anti_slave_0_address;                                             // CH3_YN1_MU_s1_translator:av_address -> CH3_YN1_MU:address
	wire          ch3_yn1_mu_s1_translator_avalon_anti_slave_0_chipselect;                                          // CH3_YN1_MU_s1_translator:av_chipselect -> CH3_YN1_MU:chipselect
	wire          ch3_yn1_mu_s1_translator_avalon_anti_slave_0_write;                                               // CH3_YN1_MU_s1_translator:av_write -> CH3_YN1_MU:write_n
	wire   [31:0] ch3_yn1_mu_s1_translator_avalon_anti_slave_0_readdata;                                            // CH3_YN1_MU:readdata -> CH3_YN1_MU_s1_translator:av_readdata
	wire   [31:0] ch3_yn1_ml_s1_translator_avalon_anti_slave_0_writedata;                                           // CH3_YN1_ML_s1_translator:av_writedata -> CH3_YN1_ML:writedata
	wire    [1:0] ch3_yn1_ml_s1_translator_avalon_anti_slave_0_address;                                             // CH3_YN1_ML_s1_translator:av_address -> CH3_YN1_ML:address
	wire          ch3_yn1_ml_s1_translator_avalon_anti_slave_0_chipselect;                                          // CH3_YN1_ML_s1_translator:av_chipselect -> CH3_YN1_ML:chipselect
	wire          ch3_yn1_ml_s1_translator_avalon_anti_slave_0_write;                                               // CH3_YN1_ML_s1_translator:av_write -> CH3_YN1_ML:write_n
	wire   [31:0] ch3_yn1_ml_s1_translator_avalon_anti_slave_0_readdata;                                            // CH3_YN1_ML:readdata -> CH3_YN1_ML_s1_translator:av_readdata
	wire   [31:0] ch4_timer_rst_s1_translator_avalon_anti_slave_0_writedata;                                        // CH4_TIMER_RST_s1_translator:av_writedata -> CH4_TIMER_RST:writedata
	wire    [1:0] ch4_timer_rst_s1_translator_avalon_anti_slave_0_address;                                          // CH4_TIMER_RST_s1_translator:av_address -> CH4_TIMER_RST:address
	wire          ch4_timer_rst_s1_translator_avalon_anti_slave_0_chipselect;                                       // CH4_TIMER_RST_s1_translator:av_chipselect -> CH4_TIMER_RST:chipselect
	wire          ch4_timer_rst_s1_translator_avalon_anti_slave_0_write;                                            // CH4_TIMER_RST_s1_translator:av_write -> CH4_TIMER_RST:write_n
	wire   [31:0] ch4_timer_rst_s1_translator_avalon_anti_slave_0_readdata;                                         // CH4_TIMER_RST:readdata -> CH4_TIMER_RST_s1_translator:av_readdata
	wire   [31:0] ch4_thresh_s1_translator_avalon_anti_slave_0_writedata;                                           // CH4_THRESH_s1_translator:av_writedata -> CH4_THRESH:writedata
	wire    [1:0] ch4_thresh_s1_translator_avalon_anti_slave_0_address;                                             // CH4_THRESH_s1_translator:av_address -> CH4_THRESH:address
	wire          ch4_thresh_s1_translator_avalon_anti_slave_0_chipselect;                                          // CH4_THRESH_s1_translator:av_chipselect -> CH4_THRESH:chipselect
	wire          ch4_thresh_s1_translator_avalon_anti_slave_0_write;                                               // CH4_THRESH_s1_translator:av_write -> CH4_THRESH:write_n
	wire   [31:0] ch4_thresh_s1_translator_avalon_anti_slave_0_readdata;                                            // CH4_THRESH:readdata -> CH4_THRESH_s1_translator:av_readdata
	wire   [31:0] ch4_rd_peak_s1_translator_avalon_anti_slave_0_writedata;                                          // CH4_RD_PEAK_s1_translator:av_writedata -> CH4_RD_PEAK:writedata
	wire    [1:0] ch4_rd_peak_s1_translator_avalon_anti_slave_0_address;                                            // CH4_RD_PEAK_s1_translator:av_address -> CH4_RD_PEAK:address
	wire          ch4_rd_peak_s1_translator_avalon_anti_slave_0_chipselect;                                         // CH4_RD_PEAK_s1_translator:av_chipselect -> CH4_RD_PEAK:chipselect
	wire          ch4_rd_peak_s1_translator_avalon_anti_slave_0_write;                                              // CH4_RD_PEAK_s1_translator:av_write -> CH4_RD_PEAK:write_n
	wire   [31:0] ch4_rd_peak_s1_translator_avalon_anti_slave_0_readdata;                                           // CH4_RD_PEAK:readdata -> CH4_RD_PEAK_s1_translator:av_readdata
	wire   [31:0] ch4_peak_found_s1_translator_avalon_anti_slave_0_writedata;                                       // CH4_PEAK_FOUND_s1_translator:av_writedata -> CH4_PEAK_FOUND:writedata
	wire    [1:0] ch4_peak_found_s1_translator_avalon_anti_slave_0_address;                                         // CH4_PEAK_FOUND_s1_translator:av_address -> CH4_PEAK_FOUND:address
	wire          ch4_peak_found_s1_translator_avalon_anti_slave_0_chipselect;                                      // CH4_PEAK_FOUND_s1_translator:av_chipselect -> CH4_PEAK_FOUND:chipselect
	wire          ch4_peak_found_s1_translator_avalon_anti_slave_0_write;                                           // CH4_PEAK_FOUND_s1_translator:av_write -> CH4_PEAK_FOUND:write_n
	wire   [31:0] ch4_peak_found_s1_translator_avalon_anti_slave_0_readdata;                                        // CH4_PEAK_FOUND:readdata -> CH4_PEAK_FOUND_s1_translator:av_readdata
	wire   [31:0] ch4_time_s1_translator_avalon_anti_slave_0_writedata;                                             // CH4_TIME_s1_translator:av_writedata -> CH4_TIME:writedata
	wire    [1:0] ch4_time_s1_translator_avalon_anti_slave_0_address;                                               // CH4_TIME_s1_translator:av_address -> CH4_TIME:address
	wire          ch4_time_s1_translator_avalon_anti_slave_0_chipselect;                                            // CH4_TIME_s1_translator:av_chipselect -> CH4_TIME:chipselect
	wire          ch4_time_s1_translator_avalon_anti_slave_0_write;                                                 // CH4_TIME_s1_translator:av_write -> CH4_TIME:write_n
	wire   [31:0] ch4_time_s1_translator_avalon_anti_slave_0_readdata;                                              // CH4_TIME:readdata -> CH4_TIME_s1_translator:av_readdata
	wire   [31:0] ch4_yn1_u_s1_translator_avalon_anti_slave_0_writedata;                                            // CH4_YN1_U_s1_translator:av_writedata -> CH4_YN1_U:writedata
	wire    [1:0] ch4_yn1_u_s1_translator_avalon_anti_slave_0_address;                                              // CH4_YN1_U_s1_translator:av_address -> CH4_YN1_U:address
	wire          ch4_yn1_u_s1_translator_avalon_anti_slave_0_chipselect;                                           // CH4_YN1_U_s1_translator:av_chipselect -> CH4_YN1_U:chipselect
	wire          ch4_yn1_u_s1_translator_avalon_anti_slave_0_write;                                                // CH4_YN1_U_s1_translator:av_write -> CH4_YN1_U:write_n
	wire   [31:0] ch4_yn1_u_s1_translator_avalon_anti_slave_0_readdata;                                             // CH4_YN1_U:readdata -> CH4_YN1_U_s1_translator:av_readdata
	wire   [31:0] ch4_yn1_mu_s1_translator_avalon_anti_slave_0_writedata;                                           // CH4_YN1_MU_s1_translator:av_writedata -> CH4_YN1_MU:writedata
	wire    [1:0] ch4_yn1_mu_s1_translator_avalon_anti_slave_0_address;                                             // CH4_YN1_MU_s1_translator:av_address -> CH4_YN1_MU:address
	wire          ch4_yn1_mu_s1_translator_avalon_anti_slave_0_chipselect;                                          // CH4_YN1_MU_s1_translator:av_chipselect -> CH4_YN1_MU:chipselect
	wire          ch4_yn1_mu_s1_translator_avalon_anti_slave_0_write;                                               // CH4_YN1_MU_s1_translator:av_write -> CH4_YN1_MU:write_n
	wire   [31:0] ch4_yn1_mu_s1_translator_avalon_anti_slave_0_readdata;                                            // CH4_YN1_MU:readdata -> CH4_YN1_MU_s1_translator:av_readdata
	wire   [31:0] ch4_yn1_ml_s1_translator_avalon_anti_slave_0_writedata;                                           // CH4_YN1_ML_s1_translator:av_writedata -> CH4_YN1_ML:writedata
	wire    [1:0] ch4_yn1_ml_s1_translator_avalon_anti_slave_0_address;                                             // CH4_YN1_ML_s1_translator:av_address -> CH4_YN1_ML:address
	wire          ch4_yn1_ml_s1_translator_avalon_anti_slave_0_chipselect;                                          // CH4_YN1_ML_s1_translator:av_chipselect -> CH4_YN1_ML:chipselect
	wire          ch4_yn1_ml_s1_translator_avalon_anti_slave_0_write;                                               // CH4_YN1_ML_s1_translator:av_write -> CH4_YN1_ML:write_n
	wire   [31:0] ch4_yn1_ml_s1_translator_avalon_anti_slave_0_readdata;                                            // CH4_YN1_ML:readdata -> CH4_YN1_ML_s1_translator:av_readdata
	wire   [31:0] ch4_yn1_l_s1_translator_avalon_anti_slave_0_writedata;                                            // CH4_YN1_L_s1_translator:av_writedata -> CH4_YN1_L:writedata
	wire    [1:0] ch4_yn1_l_s1_translator_avalon_anti_slave_0_address;                                              // CH4_YN1_L_s1_translator:av_address -> CH4_YN1_L:address
	wire          ch4_yn1_l_s1_translator_avalon_anti_slave_0_chipselect;                                           // CH4_YN1_L_s1_translator:av_chipselect -> CH4_YN1_L:chipselect
	wire          ch4_yn1_l_s1_translator_avalon_anti_slave_0_write;                                                // CH4_YN1_L_s1_translator:av_write -> CH4_YN1_L:write_n
	wire   [31:0] ch4_yn1_l_s1_translator_avalon_anti_slave_0_readdata;                                             // CH4_YN1_L:readdata -> CH4_YN1_L_s1_translator:av_readdata
	wire   [31:0] ch4_yn2_u_s1_translator_avalon_anti_slave_0_writedata;                                            // CH4_YN2_U_s1_translator:av_writedata -> CH4_YN2_U:writedata
	wire    [1:0] ch4_yn2_u_s1_translator_avalon_anti_slave_0_address;                                              // CH4_YN2_U_s1_translator:av_address -> CH4_YN2_U:address
	wire          ch4_yn2_u_s1_translator_avalon_anti_slave_0_chipselect;                                           // CH4_YN2_U_s1_translator:av_chipselect -> CH4_YN2_U:chipselect
	wire          ch4_yn2_u_s1_translator_avalon_anti_slave_0_write;                                                // CH4_YN2_U_s1_translator:av_write -> CH4_YN2_U:write_n
	wire   [31:0] ch4_yn2_u_s1_translator_avalon_anti_slave_0_readdata;                                             // CH4_YN2_U:readdata -> CH4_YN2_U_s1_translator:av_readdata
	wire   [31:0] ch4_yn2_mu_s1_translator_avalon_anti_slave_0_writedata;                                           // CH4_YN2_MU_s1_translator:av_writedata -> CH4_YN2_MU:writedata
	wire    [1:0] ch4_yn2_mu_s1_translator_avalon_anti_slave_0_address;                                             // CH4_YN2_MU_s1_translator:av_address -> CH4_YN2_MU:address
	wire          ch4_yn2_mu_s1_translator_avalon_anti_slave_0_chipselect;                                          // CH4_YN2_MU_s1_translator:av_chipselect -> CH4_YN2_MU:chipselect
	wire          ch4_yn2_mu_s1_translator_avalon_anti_slave_0_write;                                               // CH4_YN2_MU_s1_translator:av_write -> CH4_YN2_MU:write_n
	wire   [31:0] ch4_yn2_mu_s1_translator_avalon_anti_slave_0_readdata;                                            // CH4_YN2_MU:readdata -> CH4_YN2_MU_s1_translator:av_readdata
	wire   [31:0] ch4_yn2_ml_s1_translator_avalon_anti_slave_0_writedata;                                           // CH4_YN2_ML_s1_translator:av_writedata -> CH4_YN2_ML:writedata
	wire    [1:0] ch4_yn2_ml_s1_translator_avalon_anti_slave_0_address;                                             // CH4_YN2_ML_s1_translator:av_address -> CH4_YN2_ML:address
	wire          ch4_yn2_ml_s1_translator_avalon_anti_slave_0_chipselect;                                          // CH4_YN2_ML_s1_translator:av_chipselect -> CH4_YN2_ML:chipselect
	wire          ch4_yn2_ml_s1_translator_avalon_anti_slave_0_write;                                               // CH4_YN2_ML_s1_translator:av_write -> CH4_YN2_ML:write_n
	wire   [31:0] ch4_yn2_ml_s1_translator_avalon_anti_slave_0_readdata;                                            // CH4_YN2_ML:readdata -> CH4_YN2_ML_s1_translator:av_readdata
	wire   [31:0] ch4_yn2_l_s1_translator_avalon_anti_slave_0_writedata;                                            // CH4_YN2_L_s1_translator:av_writedata -> CH4_YN2_L:writedata
	wire    [1:0] ch4_yn2_l_s1_translator_avalon_anti_slave_0_address;                                              // CH4_YN2_L_s1_translator:av_address -> CH4_YN2_L:address
	wire          ch4_yn2_l_s1_translator_avalon_anti_slave_0_chipselect;                                           // CH4_YN2_L_s1_translator:av_chipselect -> CH4_YN2_L:chipselect
	wire          ch4_yn2_l_s1_translator_avalon_anti_slave_0_write;                                                // CH4_YN2_L_s1_translator:av_write -> CH4_YN2_L:write_n
	wire   [31:0] ch4_yn2_l_s1_translator_avalon_anti_slave_0_readdata;                                             // CH4_YN2_L:readdata -> CH4_YN2_L_s1_translator:av_readdata
	wire   [31:0] ch4_yn3_u_s1_translator_avalon_anti_slave_0_writedata;                                            // CH4_YN3_U_s1_translator:av_writedata -> CH4_YN3_U:writedata
	wire    [1:0] ch4_yn3_u_s1_translator_avalon_anti_slave_0_address;                                              // CH4_YN3_U_s1_translator:av_address -> CH4_YN3_U:address
	wire          ch4_yn3_u_s1_translator_avalon_anti_slave_0_chipselect;                                           // CH4_YN3_U_s1_translator:av_chipselect -> CH4_YN3_U:chipselect
	wire          ch4_yn3_u_s1_translator_avalon_anti_slave_0_write;                                                // CH4_YN3_U_s1_translator:av_write -> CH4_YN3_U:write_n
	wire   [31:0] ch4_yn3_u_s1_translator_avalon_anti_slave_0_readdata;                                             // CH4_YN3_U:readdata -> CH4_YN3_U_s1_translator:av_readdata
	wire   [31:0] ch4_yn3_mu_s1_translator_avalon_anti_slave_0_writedata;                                           // CH4_YN3_MU_s1_translator:av_writedata -> CH4_YN3_MU:writedata
	wire    [1:0] ch4_yn3_mu_s1_translator_avalon_anti_slave_0_address;                                             // CH4_YN3_MU_s1_translator:av_address -> CH4_YN3_MU:address
	wire          ch4_yn3_mu_s1_translator_avalon_anti_slave_0_chipselect;                                          // CH4_YN3_MU_s1_translator:av_chipselect -> CH4_YN3_MU:chipselect
	wire          ch4_yn3_mu_s1_translator_avalon_anti_slave_0_write;                                               // CH4_YN3_MU_s1_translator:av_write -> CH4_YN3_MU:write_n
	wire   [31:0] ch4_yn3_mu_s1_translator_avalon_anti_slave_0_readdata;                                            // CH4_YN3_MU:readdata -> CH4_YN3_MU_s1_translator:av_readdata
	wire   [31:0] ch4_yn3_ml_s1_translator_avalon_anti_slave_0_writedata;                                           // CH4_YN3_ML_s1_translator:av_writedata -> CH4_YN3_ML:writedata
	wire    [1:0] ch4_yn3_ml_s1_translator_avalon_anti_slave_0_address;                                             // CH4_YN3_ML_s1_translator:av_address -> CH4_YN3_ML:address
	wire          ch4_yn3_ml_s1_translator_avalon_anti_slave_0_chipselect;                                          // CH4_YN3_ML_s1_translator:av_chipselect -> CH4_YN3_ML:chipselect
	wire          ch4_yn3_ml_s1_translator_avalon_anti_slave_0_write;                                               // CH4_YN3_ML_s1_translator:av_write -> CH4_YN3_ML:write_n
	wire   [31:0] ch4_yn3_ml_s1_translator_avalon_anti_slave_0_readdata;                                            // CH4_YN3_ML:readdata -> CH4_YN3_ML_s1_translator:av_readdata
	wire   [31:0] ch4_yn3_l_s1_translator_avalon_anti_slave_0_writedata;                                            // CH4_YN3_L_s1_translator:av_writedata -> CH4_YN3_L:writedata
	wire    [1:0] ch4_yn3_l_s1_translator_avalon_anti_slave_0_address;                                              // CH4_YN3_L_s1_translator:av_address -> CH4_YN3_L:address
	wire          ch4_yn3_l_s1_translator_avalon_anti_slave_0_chipselect;                                           // CH4_YN3_L_s1_translator:av_chipselect -> CH4_YN3_L:chipselect
	wire          ch4_yn3_l_s1_translator_avalon_anti_slave_0_write;                                                // CH4_YN3_L_s1_translator:av_write -> CH4_YN3_L:write_n
	wire   [31:0] ch4_yn3_l_s1_translator_avalon_anti_slave_0_readdata;                                             // CH4_YN3_L:readdata -> CH4_YN3_L_s1_translator:av_readdata
	wire          nios_cpu_instruction_master_translator_avalon_universal_master_0_waitrequest;                     // NIOS_CPU_instruction_master_translator_avalon_universal_master_0_agent:av_waitrequest -> NIOS_CPU_instruction_master_translator:uav_waitrequest
	wire    [2:0] nios_cpu_instruction_master_translator_avalon_universal_master_0_burstcount;                      // NIOS_CPU_instruction_master_translator:uav_burstcount -> NIOS_CPU_instruction_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] nios_cpu_instruction_master_translator_avalon_universal_master_0_writedata;                       // NIOS_CPU_instruction_master_translator:uav_writedata -> NIOS_CPU_instruction_master_translator_avalon_universal_master_0_agent:av_writedata
	wire   [21:0] nios_cpu_instruction_master_translator_avalon_universal_master_0_address;                         // NIOS_CPU_instruction_master_translator:uav_address -> NIOS_CPU_instruction_master_translator_avalon_universal_master_0_agent:av_address
	wire          nios_cpu_instruction_master_translator_avalon_universal_master_0_lock;                            // NIOS_CPU_instruction_master_translator:uav_lock -> NIOS_CPU_instruction_master_translator_avalon_universal_master_0_agent:av_lock
	wire          nios_cpu_instruction_master_translator_avalon_universal_master_0_write;                           // NIOS_CPU_instruction_master_translator:uav_write -> NIOS_CPU_instruction_master_translator_avalon_universal_master_0_agent:av_write
	wire          nios_cpu_instruction_master_translator_avalon_universal_master_0_read;                            // NIOS_CPU_instruction_master_translator:uav_read -> NIOS_CPU_instruction_master_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] nios_cpu_instruction_master_translator_avalon_universal_master_0_readdata;                        // NIOS_CPU_instruction_master_translator_avalon_universal_master_0_agent:av_readdata -> NIOS_CPU_instruction_master_translator:uav_readdata
	wire          nios_cpu_instruction_master_translator_avalon_universal_master_0_debugaccess;                     // NIOS_CPU_instruction_master_translator:uav_debugaccess -> NIOS_CPU_instruction_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] nios_cpu_instruction_master_translator_avalon_universal_master_0_byteenable;                      // NIOS_CPU_instruction_master_translator:uav_byteenable -> NIOS_CPU_instruction_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire          nios_cpu_instruction_master_translator_avalon_universal_master_0_readdatavalid;                   // NIOS_CPU_instruction_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> NIOS_CPU_instruction_master_translator:uav_readdatavalid
	wire          nios_cpu_data_master_translator_avalon_universal_master_0_waitrequest;                            // NIOS_CPU_data_master_translator_avalon_universal_master_0_agent:av_waitrequest -> NIOS_CPU_data_master_translator:uav_waitrequest
	wire    [2:0] nios_cpu_data_master_translator_avalon_universal_master_0_burstcount;                             // NIOS_CPU_data_master_translator:uav_burstcount -> NIOS_CPU_data_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] nios_cpu_data_master_translator_avalon_universal_master_0_writedata;                              // NIOS_CPU_data_master_translator:uav_writedata -> NIOS_CPU_data_master_translator_avalon_universal_master_0_agent:av_writedata
	wire   [21:0] nios_cpu_data_master_translator_avalon_universal_master_0_address;                                // NIOS_CPU_data_master_translator:uav_address -> NIOS_CPU_data_master_translator_avalon_universal_master_0_agent:av_address
	wire          nios_cpu_data_master_translator_avalon_universal_master_0_lock;                                   // NIOS_CPU_data_master_translator:uav_lock -> NIOS_CPU_data_master_translator_avalon_universal_master_0_agent:av_lock
	wire          nios_cpu_data_master_translator_avalon_universal_master_0_write;                                  // NIOS_CPU_data_master_translator:uav_write -> NIOS_CPU_data_master_translator_avalon_universal_master_0_agent:av_write
	wire          nios_cpu_data_master_translator_avalon_universal_master_0_read;                                   // NIOS_CPU_data_master_translator:uav_read -> NIOS_CPU_data_master_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] nios_cpu_data_master_translator_avalon_universal_master_0_readdata;                               // NIOS_CPU_data_master_translator_avalon_universal_master_0_agent:av_readdata -> NIOS_CPU_data_master_translator:uav_readdata
	wire          nios_cpu_data_master_translator_avalon_universal_master_0_debugaccess;                            // NIOS_CPU_data_master_translator:uav_debugaccess -> NIOS_CPU_data_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] nios_cpu_data_master_translator_avalon_universal_master_0_byteenable;                             // NIOS_CPU_data_master_translator:uav_byteenable -> NIOS_CPU_data_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire          nios_cpu_data_master_translator_avalon_universal_master_0_readdatavalid;                          // NIOS_CPU_data_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> NIOS_CPU_data_master_translator:uav_readdatavalid
	wire          nios_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest;              // NIOS_CPU_jtag_debug_module_translator:uav_waitrequest -> NIOS_CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] nios_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount;               // NIOS_CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_burstcount -> NIOS_CPU_jtag_debug_module_translator:uav_burstcount
	wire   [31:0] nios_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata;                // NIOS_CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_writedata -> NIOS_CPU_jtag_debug_module_translator:uav_writedata
	wire   [21:0] nios_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address;                  // NIOS_CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_address -> NIOS_CPU_jtag_debug_module_translator:uav_address
	wire          nios_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write;                    // NIOS_CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_write -> NIOS_CPU_jtag_debug_module_translator:uav_write
	wire          nios_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock;                     // NIOS_CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_lock -> NIOS_CPU_jtag_debug_module_translator:uav_lock
	wire          nios_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read;                     // NIOS_CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_read -> NIOS_CPU_jtag_debug_module_translator:uav_read
	wire   [31:0] nios_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata;                 // NIOS_CPU_jtag_debug_module_translator:uav_readdata -> NIOS_CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          nios_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid;            // NIOS_CPU_jtag_debug_module_translator:uav_readdatavalid -> NIOS_CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          nios_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess;              // NIOS_CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_debugaccess -> NIOS_CPU_jtag_debug_module_translator:uav_debugaccess
	wire    [3:0] nios_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable;               // NIOS_CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_byteenable -> NIOS_CPU_jtag_debug_module_translator:uav_byteenable
	wire          nios_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;       // NIOS_CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> NIOS_CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          nios_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid;             // NIOS_CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_valid -> NIOS_CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          nios_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;     // NIOS_CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> NIOS_CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] nios_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data;              // NIOS_CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_data -> NIOS_CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          nios_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready;             // NIOS_CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> NIOS_CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          nios_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;    // NIOS_CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> NIOS_CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          nios_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;          // NIOS_CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> NIOS_CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          nios_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;  // NIOS_CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> NIOS_CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] nios_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;           // NIOS_CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> NIOS_CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          nios_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;          // NIOS_CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_ready -> NIOS_CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          nios_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;        // NIOS_CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> NIOS_CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] nios_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;         // NIOS_CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> NIOS_CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          nios_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;        // NIOS_CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> NIOS_CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          ram_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                  // RAM_s1_translator:uav_waitrequest -> RAM_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] ram_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                   // RAM_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> RAM_s1_translator:uav_burstcount
	wire   [31:0] ram_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                    // RAM_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> RAM_s1_translator:uav_writedata
	wire   [21:0] ram_s1_translator_avalon_universal_slave_0_agent_m0_address;                                      // RAM_s1_translator_avalon_universal_slave_0_agent:m0_address -> RAM_s1_translator:uav_address
	wire          ram_s1_translator_avalon_universal_slave_0_agent_m0_write;                                        // RAM_s1_translator_avalon_universal_slave_0_agent:m0_write -> RAM_s1_translator:uav_write
	wire          ram_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                         // RAM_s1_translator_avalon_universal_slave_0_agent:m0_lock -> RAM_s1_translator:uav_lock
	wire          ram_s1_translator_avalon_universal_slave_0_agent_m0_read;                                         // RAM_s1_translator_avalon_universal_slave_0_agent:m0_read -> RAM_s1_translator:uav_read
	wire   [31:0] ram_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                     // RAM_s1_translator:uav_readdata -> RAM_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          ram_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                // RAM_s1_translator:uav_readdatavalid -> RAM_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          ram_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                  // RAM_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> RAM_s1_translator:uav_debugaccess
	wire    [3:0] ram_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                   // RAM_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> RAM_s1_translator:uav_byteenable
	wire          ram_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                           // RAM_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> RAM_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          ram_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                 // RAM_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> RAM_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          ram_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                         // RAM_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> RAM_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] ram_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                  // RAM_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> RAM_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          ram_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                 // RAM_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> RAM_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                        // RAM_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> RAM_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                              // RAM_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> RAM_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                      // RAM_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> RAM_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                               // RAM_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> RAM_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                              // RAM_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> RAM_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          ram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                            // RAM_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> RAM_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] ram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                             // RAM_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> RAM_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          ram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                            // RAM_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> RAM_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          ssram_uas_translator_avalon_universal_slave_0_agent_m0_waitrequest;                               // SSRAM_uas_translator:uav_waitrequest -> SSRAM_uas_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] ssram_uas_translator_avalon_universal_slave_0_agent_m0_burstcount;                                // SSRAM_uas_translator_avalon_universal_slave_0_agent:m0_burstcount -> SSRAM_uas_translator:uav_burstcount
	wire   [31:0] ssram_uas_translator_avalon_universal_slave_0_agent_m0_writedata;                                 // SSRAM_uas_translator_avalon_universal_slave_0_agent:m0_writedata -> SSRAM_uas_translator:uav_writedata
	wire   [21:0] ssram_uas_translator_avalon_universal_slave_0_agent_m0_address;                                   // SSRAM_uas_translator_avalon_universal_slave_0_agent:m0_address -> SSRAM_uas_translator:uav_address
	wire          ssram_uas_translator_avalon_universal_slave_0_agent_m0_write;                                     // SSRAM_uas_translator_avalon_universal_slave_0_agent:m0_write -> SSRAM_uas_translator:uav_write
	wire          ssram_uas_translator_avalon_universal_slave_0_agent_m0_lock;                                      // SSRAM_uas_translator_avalon_universal_slave_0_agent:m0_lock -> SSRAM_uas_translator:uav_lock
	wire          ssram_uas_translator_avalon_universal_slave_0_agent_m0_read;                                      // SSRAM_uas_translator_avalon_universal_slave_0_agent:m0_read -> SSRAM_uas_translator:uav_read
	wire   [31:0] ssram_uas_translator_avalon_universal_slave_0_agent_m0_readdata;                                  // SSRAM_uas_translator:uav_readdata -> SSRAM_uas_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          ssram_uas_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                             // SSRAM_uas_translator:uav_readdatavalid -> SSRAM_uas_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          ssram_uas_translator_avalon_universal_slave_0_agent_m0_debugaccess;                               // SSRAM_uas_translator_avalon_universal_slave_0_agent:m0_debugaccess -> SSRAM_uas_translator:uav_debugaccess
	wire    [3:0] ssram_uas_translator_avalon_universal_slave_0_agent_m0_byteenable;                                // SSRAM_uas_translator_avalon_universal_slave_0_agent:m0_byteenable -> SSRAM_uas_translator:uav_byteenable
	wire          ssram_uas_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                        // SSRAM_uas_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> SSRAM_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          ssram_uas_translator_avalon_universal_slave_0_agent_rf_source_valid;                              // SSRAM_uas_translator_avalon_universal_slave_0_agent:rf_source_valid -> SSRAM_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          ssram_uas_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                      // SSRAM_uas_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> SSRAM_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] ssram_uas_translator_avalon_universal_slave_0_agent_rf_source_data;                               // SSRAM_uas_translator_avalon_universal_slave_0_agent:rf_source_data -> SSRAM_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          ssram_uas_translator_avalon_universal_slave_0_agent_rf_source_ready;                              // SSRAM_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> SSRAM_uas_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          ssram_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                     // SSRAM_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> SSRAM_uas_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          ssram_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                           // SSRAM_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> SSRAM_uas_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          ssram_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                   // SSRAM_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> SSRAM_uas_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] ssram_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                            // SSRAM_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> SSRAM_uas_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          ssram_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                           // SSRAM_uas_translator_avalon_universal_slave_0_agent:rf_sink_ready -> SSRAM_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          ssram_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                         // SSRAM_uas_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> SSRAM_uas_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] ssram_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                          // SSRAM_uas_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> SSRAM_uas_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          ssram_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                         // SSRAM_uas_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> SSRAM_uas_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;             // JTAG_UART_avalon_jtag_slave_translator:uav_waitrequest -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;              // JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> JTAG_UART_avalon_jtag_slave_translator:uav_burstcount
	wire   [31:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata;               // JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> JTAG_UART_avalon_jtag_slave_translator:uav_writedata
	wire   [21:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address;                 // JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_address -> JTAG_UART_avalon_jtag_slave_translator:uav_address
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write;                   // JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_write -> JTAG_UART_avalon_jtag_slave_translator:uav_write
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock;                    // JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_lock -> JTAG_UART_avalon_jtag_slave_translator:uav_lock
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read;                    // JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_read -> JTAG_UART_avalon_jtag_slave_translator:uav_read
	wire   [31:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                // JTAG_UART_avalon_jtag_slave_translator:uav_readdata -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;           // JTAG_UART_avalon_jtag_slave_translator:uav_readdatavalid -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;             // JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> JTAG_UART_avalon_jtag_slave_translator:uav_debugaccess
	wire    [3:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;              // JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> JTAG_UART_avalon_jtag_slave_translator:uav_byteenable
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;      // JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;            // JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;    // JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data;             // JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;            // JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;   // JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;         // JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket; // JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;          // JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;         // JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;       // JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;        // JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;       // JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                       // LCD_control_slave_translator:uav_waitrequest -> LCD_control_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                        // LCD_control_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> LCD_control_slave_translator:uav_burstcount
	wire   [31:0] lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                         // LCD_control_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> LCD_control_slave_translator:uav_writedata
	wire   [21:0] lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_address;                           // LCD_control_slave_translator_avalon_universal_slave_0_agent:m0_address -> LCD_control_slave_translator:uav_address
	wire          lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_write;                             // LCD_control_slave_translator_avalon_universal_slave_0_agent:m0_write -> LCD_control_slave_translator:uav_write
	wire          lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_lock;                              // LCD_control_slave_translator_avalon_universal_slave_0_agent:m0_lock -> LCD_control_slave_translator:uav_lock
	wire          lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_read;                              // LCD_control_slave_translator_avalon_universal_slave_0_agent:m0_read -> LCD_control_slave_translator:uav_read
	wire   [31:0] lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                          // LCD_control_slave_translator:uav_readdata -> LCD_control_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                     // LCD_control_slave_translator:uav_readdatavalid -> LCD_control_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                       // LCD_control_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> LCD_control_slave_translator:uav_debugaccess
	wire    [3:0] lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                        // LCD_control_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> LCD_control_slave_translator:uav_byteenable
	wire          lcd_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                // LCD_control_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> LCD_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          lcd_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                      // LCD_control_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> LCD_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          lcd_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;              // LCD_control_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> LCD_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] lcd_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                       // LCD_control_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> LCD_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          lcd_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                      // LCD_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> LCD_control_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;             // LCD_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> LCD_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                   // LCD_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> LCD_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;           // LCD_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> LCD_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                    // LCD_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> LCD_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                   // LCD_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> LCD_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          lcd_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                 // LCD_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> LCD_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] lcd_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                  // LCD_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> LCD_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          lcd_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                 // LCD_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> LCD_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          adc_on_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                               // ADC_ON_s1_translator:uav_waitrequest -> ADC_ON_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] adc_on_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                // ADC_ON_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> ADC_ON_s1_translator:uav_burstcount
	wire   [31:0] adc_on_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                 // ADC_ON_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> ADC_ON_s1_translator:uav_writedata
	wire   [21:0] adc_on_s1_translator_avalon_universal_slave_0_agent_m0_address;                                   // ADC_ON_s1_translator_avalon_universal_slave_0_agent:m0_address -> ADC_ON_s1_translator:uav_address
	wire          adc_on_s1_translator_avalon_universal_slave_0_agent_m0_write;                                     // ADC_ON_s1_translator_avalon_universal_slave_0_agent:m0_write -> ADC_ON_s1_translator:uav_write
	wire          adc_on_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                      // ADC_ON_s1_translator_avalon_universal_slave_0_agent:m0_lock -> ADC_ON_s1_translator:uav_lock
	wire          adc_on_s1_translator_avalon_universal_slave_0_agent_m0_read;                                      // ADC_ON_s1_translator_avalon_universal_slave_0_agent:m0_read -> ADC_ON_s1_translator:uav_read
	wire   [31:0] adc_on_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                  // ADC_ON_s1_translator:uav_readdata -> ADC_ON_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          adc_on_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                             // ADC_ON_s1_translator:uav_readdatavalid -> ADC_ON_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          adc_on_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                               // ADC_ON_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> ADC_ON_s1_translator:uav_debugaccess
	wire    [3:0] adc_on_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                // ADC_ON_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> ADC_ON_s1_translator:uav_byteenable
	wire          adc_on_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                        // ADC_ON_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> ADC_ON_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          adc_on_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                              // ADC_ON_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> ADC_ON_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          adc_on_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                      // ADC_ON_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> ADC_ON_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] adc_on_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                               // ADC_ON_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> ADC_ON_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          adc_on_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                              // ADC_ON_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> ADC_ON_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          adc_on_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                     // ADC_ON_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> ADC_ON_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          adc_on_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                           // ADC_ON_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> ADC_ON_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          adc_on_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                   // ADC_ON_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> ADC_ON_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] adc_on_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                            // ADC_ON_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> ADC_ON_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          adc_on_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                           // ADC_ON_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> ADC_ON_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          adc_on_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                         // ADC_ON_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> ADC_ON_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] adc_on_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                          // ADC_ON_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> ADC_ON_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          adc_on_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                         // ADC_ON_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> ADC_ON_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          fifo_adc_data_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                        // FIFO_ADC_DATA_s1_translator:uav_waitrequest -> FIFO_ADC_DATA_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] fifo_adc_data_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                         // FIFO_ADC_DATA_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> FIFO_ADC_DATA_s1_translator:uav_burstcount
	wire   [31:0] fifo_adc_data_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                          // FIFO_ADC_DATA_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> FIFO_ADC_DATA_s1_translator:uav_writedata
	wire   [21:0] fifo_adc_data_s1_translator_avalon_universal_slave_0_agent_m0_address;                            // FIFO_ADC_DATA_s1_translator_avalon_universal_slave_0_agent:m0_address -> FIFO_ADC_DATA_s1_translator:uav_address
	wire          fifo_adc_data_s1_translator_avalon_universal_slave_0_agent_m0_write;                              // FIFO_ADC_DATA_s1_translator_avalon_universal_slave_0_agent:m0_write -> FIFO_ADC_DATA_s1_translator:uav_write
	wire          fifo_adc_data_s1_translator_avalon_universal_slave_0_agent_m0_lock;                               // FIFO_ADC_DATA_s1_translator_avalon_universal_slave_0_agent:m0_lock -> FIFO_ADC_DATA_s1_translator:uav_lock
	wire          fifo_adc_data_s1_translator_avalon_universal_slave_0_agent_m0_read;                               // FIFO_ADC_DATA_s1_translator_avalon_universal_slave_0_agent:m0_read -> FIFO_ADC_DATA_s1_translator:uav_read
	wire   [31:0] fifo_adc_data_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                           // FIFO_ADC_DATA_s1_translator:uav_readdata -> FIFO_ADC_DATA_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          fifo_adc_data_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                      // FIFO_ADC_DATA_s1_translator:uav_readdatavalid -> FIFO_ADC_DATA_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          fifo_adc_data_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                        // FIFO_ADC_DATA_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> FIFO_ADC_DATA_s1_translator:uav_debugaccess
	wire    [3:0] fifo_adc_data_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                         // FIFO_ADC_DATA_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> FIFO_ADC_DATA_s1_translator:uav_byteenable
	wire          fifo_adc_data_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                 // FIFO_ADC_DATA_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> FIFO_ADC_DATA_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          fifo_adc_data_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                       // FIFO_ADC_DATA_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> FIFO_ADC_DATA_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          fifo_adc_data_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;               // FIFO_ADC_DATA_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> FIFO_ADC_DATA_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] fifo_adc_data_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                        // FIFO_ADC_DATA_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> FIFO_ADC_DATA_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          fifo_adc_data_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                       // FIFO_ADC_DATA_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> FIFO_ADC_DATA_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          fifo_adc_data_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;              // FIFO_ADC_DATA_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> FIFO_ADC_DATA_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          fifo_adc_data_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                    // FIFO_ADC_DATA_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> FIFO_ADC_DATA_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          fifo_adc_data_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;            // FIFO_ADC_DATA_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> FIFO_ADC_DATA_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] fifo_adc_data_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                     // FIFO_ADC_DATA_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> FIFO_ADC_DATA_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          fifo_adc_data_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                    // FIFO_ADC_DATA_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> FIFO_ADC_DATA_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          fifo_adc_data_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                  // FIFO_ADC_DATA_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> FIFO_ADC_DATA_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] fifo_adc_data_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                   // FIFO_ADC_DATA_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> FIFO_ADC_DATA_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          fifo_adc_data_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                  // FIFO_ADC_DATA_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> FIFO_ADC_DATA_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          fifo_adc_data_valid_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                  // FIFO_ADC_DATA_VALID_s1_translator:uav_waitrequest -> FIFO_ADC_DATA_VALID_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] fifo_adc_data_valid_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                   // FIFO_ADC_DATA_VALID_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> FIFO_ADC_DATA_VALID_s1_translator:uav_burstcount
	wire   [31:0] fifo_adc_data_valid_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                    // FIFO_ADC_DATA_VALID_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> FIFO_ADC_DATA_VALID_s1_translator:uav_writedata
	wire   [21:0] fifo_adc_data_valid_s1_translator_avalon_universal_slave_0_agent_m0_address;                      // FIFO_ADC_DATA_VALID_s1_translator_avalon_universal_slave_0_agent:m0_address -> FIFO_ADC_DATA_VALID_s1_translator:uav_address
	wire          fifo_adc_data_valid_s1_translator_avalon_universal_slave_0_agent_m0_write;                        // FIFO_ADC_DATA_VALID_s1_translator_avalon_universal_slave_0_agent:m0_write -> FIFO_ADC_DATA_VALID_s1_translator:uav_write
	wire          fifo_adc_data_valid_s1_translator_avalon_universal_slave_0_agent_m0_lock;                         // FIFO_ADC_DATA_VALID_s1_translator_avalon_universal_slave_0_agent:m0_lock -> FIFO_ADC_DATA_VALID_s1_translator:uav_lock
	wire          fifo_adc_data_valid_s1_translator_avalon_universal_slave_0_agent_m0_read;                         // FIFO_ADC_DATA_VALID_s1_translator_avalon_universal_slave_0_agent:m0_read -> FIFO_ADC_DATA_VALID_s1_translator:uav_read
	wire   [31:0] fifo_adc_data_valid_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                     // FIFO_ADC_DATA_VALID_s1_translator:uav_readdata -> FIFO_ADC_DATA_VALID_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          fifo_adc_data_valid_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                // FIFO_ADC_DATA_VALID_s1_translator:uav_readdatavalid -> FIFO_ADC_DATA_VALID_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          fifo_adc_data_valid_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                  // FIFO_ADC_DATA_VALID_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> FIFO_ADC_DATA_VALID_s1_translator:uav_debugaccess
	wire    [3:0] fifo_adc_data_valid_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                   // FIFO_ADC_DATA_VALID_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> FIFO_ADC_DATA_VALID_s1_translator:uav_byteenable
	wire          fifo_adc_data_valid_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;           // FIFO_ADC_DATA_VALID_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> FIFO_ADC_DATA_VALID_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          fifo_adc_data_valid_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                 // FIFO_ADC_DATA_VALID_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> FIFO_ADC_DATA_VALID_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          fifo_adc_data_valid_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;         // FIFO_ADC_DATA_VALID_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> FIFO_ADC_DATA_VALID_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] fifo_adc_data_valid_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                  // FIFO_ADC_DATA_VALID_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> FIFO_ADC_DATA_VALID_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          fifo_adc_data_valid_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                 // FIFO_ADC_DATA_VALID_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> FIFO_ADC_DATA_VALID_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          fifo_adc_data_valid_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;        // FIFO_ADC_DATA_VALID_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> FIFO_ADC_DATA_VALID_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          fifo_adc_data_valid_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;              // FIFO_ADC_DATA_VALID_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> FIFO_ADC_DATA_VALID_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          fifo_adc_data_valid_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;      // FIFO_ADC_DATA_VALID_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> FIFO_ADC_DATA_VALID_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] fifo_adc_data_valid_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;               // FIFO_ADC_DATA_VALID_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> FIFO_ADC_DATA_VALID_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          fifo_adc_data_valid_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;              // FIFO_ADC_DATA_VALID_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> FIFO_ADC_DATA_VALID_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          fifo_adc_data_valid_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;            // FIFO_ADC_DATA_VALID_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> FIFO_ADC_DATA_VALID_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] fifo_adc_data_valid_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;             // FIFO_ADC_DATA_VALID_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> FIFO_ADC_DATA_VALID_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          fifo_adc_data_valid_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;            // FIFO_ADC_DATA_VALID_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> FIFO_ADC_DATA_VALID_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          fifo_rst_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                             // FIFO_RST_s1_translator:uav_waitrequest -> FIFO_RST_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] fifo_rst_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                              // FIFO_RST_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> FIFO_RST_s1_translator:uav_burstcount
	wire   [31:0] fifo_rst_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                               // FIFO_RST_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> FIFO_RST_s1_translator:uav_writedata
	wire   [21:0] fifo_rst_s1_translator_avalon_universal_slave_0_agent_m0_address;                                 // FIFO_RST_s1_translator_avalon_universal_slave_0_agent:m0_address -> FIFO_RST_s1_translator:uav_address
	wire          fifo_rst_s1_translator_avalon_universal_slave_0_agent_m0_write;                                   // FIFO_RST_s1_translator_avalon_universal_slave_0_agent:m0_write -> FIFO_RST_s1_translator:uav_write
	wire          fifo_rst_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                    // FIFO_RST_s1_translator_avalon_universal_slave_0_agent:m0_lock -> FIFO_RST_s1_translator:uav_lock
	wire          fifo_rst_s1_translator_avalon_universal_slave_0_agent_m0_read;                                    // FIFO_RST_s1_translator_avalon_universal_slave_0_agent:m0_read -> FIFO_RST_s1_translator:uav_read
	wire   [31:0] fifo_rst_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                // FIFO_RST_s1_translator:uav_readdata -> FIFO_RST_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          fifo_rst_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                           // FIFO_RST_s1_translator:uav_readdatavalid -> FIFO_RST_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          fifo_rst_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                             // FIFO_RST_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> FIFO_RST_s1_translator:uav_debugaccess
	wire    [3:0] fifo_rst_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                              // FIFO_RST_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> FIFO_RST_s1_translator:uav_byteenable
	wire          fifo_rst_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                      // FIFO_RST_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> FIFO_RST_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          fifo_rst_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                            // FIFO_RST_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> FIFO_RST_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          fifo_rst_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                    // FIFO_RST_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> FIFO_RST_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] fifo_rst_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                             // FIFO_RST_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> FIFO_RST_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          fifo_rst_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                            // FIFO_RST_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> FIFO_RST_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          fifo_rst_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                   // FIFO_RST_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> FIFO_RST_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          fifo_rst_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                         // FIFO_RST_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> FIFO_RST_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          fifo_rst_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                 // FIFO_RST_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> FIFO_RST_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] fifo_rst_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                          // FIFO_RST_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> FIFO_RST_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          fifo_rst_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                         // FIFO_RST_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> FIFO_RST_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          fifo_rst_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                       // FIFO_RST_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> FIFO_RST_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] fifo_rst_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                        // FIFO_RST_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> FIFO_RST_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          fifo_rst_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                       // FIFO_RST_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> FIFO_RST_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          subtractor_on_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                        // SUBTRACTOR_ON_s1_translator:uav_waitrequest -> SUBTRACTOR_ON_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] subtractor_on_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                         // SUBTRACTOR_ON_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> SUBTRACTOR_ON_s1_translator:uav_burstcount
	wire   [31:0] subtractor_on_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                          // SUBTRACTOR_ON_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> SUBTRACTOR_ON_s1_translator:uav_writedata
	wire   [21:0] subtractor_on_s1_translator_avalon_universal_slave_0_agent_m0_address;                            // SUBTRACTOR_ON_s1_translator_avalon_universal_slave_0_agent:m0_address -> SUBTRACTOR_ON_s1_translator:uav_address
	wire          subtractor_on_s1_translator_avalon_universal_slave_0_agent_m0_write;                              // SUBTRACTOR_ON_s1_translator_avalon_universal_slave_0_agent:m0_write -> SUBTRACTOR_ON_s1_translator:uav_write
	wire          subtractor_on_s1_translator_avalon_universal_slave_0_agent_m0_lock;                               // SUBTRACTOR_ON_s1_translator_avalon_universal_slave_0_agent:m0_lock -> SUBTRACTOR_ON_s1_translator:uav_lock
	wire          subtractor_on_s1_translator_avalon_universal_slave_0_agent_m0_read;                               // SUBTRACTOR_ON_s1_translator_avalon_universal_slave_0_agent:m0_read -> SUBTRACTOR_ON_s1_translator:uav_read
	wire   [31:0] subtractor_on_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                           // SUBTRACTOR_ON_s1_translator:uav_readdata -> SUBTRACTOR_ON_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          subtractor_on_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                      // SUBTRACTOR_ON_s1_translator:uav_readdatavalid -> SUBTRACTOR_ON_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          subtractor_on_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                        // SUBTRACTOR_ON_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> SUBTRACTOR_ON_s1_translator:uav_debugaccess
	wire    [3:0] subtractor_on_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                         // SUBTRACTOR_ON_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> SUBTRACTOR_ON_s1_translator:uav_byteenable
	wire          subtractor_on_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                 // SUBTRACTOR_ON_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> SUBTRACTOR_ON_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          subtractor_on_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                       // SUBTRACTOR_ON_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> SUBTRACTOR_ON_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          subtractor_on_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;               // SUBTRACTOR_ON_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> SUBTRACTOR_ON_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] subtractor_on_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                        // SUBTRACTOR_ON_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> SUBTRACTOR_ON_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          subtractor_on_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                       // SUBTRACTOR_ON_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> SUBTRACTOR_ON_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          subtractor_on_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;              // SUBTRACTOR_ON_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> SUBTRACTOR_ON_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          subtractor_on_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                    // SUBTRACTOR_ON_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> SUBTRACTOR_ON_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          subtractor_on_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;            // SUBTRACTOR_ON_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> SUBTRACTOR_ON_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] subtractor_on_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                     // SUBTRACTOR_ON_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> SUBTRACTOR_ON_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          subtractor_on_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                    // SUBTRACTOR_ON_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> SUBTRACTOR_ON_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          subtractor_on_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                  // SUBTRACTOR_ON_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> SUBTRACTOR_ON_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] subtractor_on_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                   // SUBTRACTOR_ON_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> SUBTRACTOR_ON_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          subtractor_on_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                  // SUBTRACTOR_ON_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> SUBTRACTOR_ON_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          ch0_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                        // CH0_TIMER_RST_s1_translator:uav_waitrequest -> CH0_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] ch0_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                         // CH0_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> CH0_TIMER_RST_s1_translator:uav_burstcount
	wire   [31:0] ch0_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                          // CH0_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> CH0_TIMER_RST_s1_translator:uav_writedata
	wire   [21:0] ch0_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_address;                            // CH0_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:m0_address -> CH0_TIMER_RST_s1_translator:uav_address
	wire          ch0_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_write;                              // CH0_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:m0_write -> CH0_TIMER_RST_s1_translator:uav_write
	wire          ch0_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_lock;                               // CH0_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:m0_lock -> CH0_TIMER_RST_s1_translator:uav_lock
	wire          ch0_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_read;                               // CH0_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:m0_read -> CH0_TIMER_RST_s1_translator:uav_read
	wire   [31:0] ch0_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                           // CH0_TIMER_RST_s1_translator:uav_readdata -> CH0_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          ch0_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                      // CH0_TIMER_RST_s1_translator:uav_readdatavalid -> CH0_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          ch0_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                        // CH0_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> CH0_TIMER_RST_s1_translator:uav_debugaccess
	wire    [3:0] ch0_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                         // CH0_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> CH0_TIMER_RST_s1_translator:uav_byteenable
	wire          ch0_timer_rst_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                 // CH0_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> CH0_TIMER_RST_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          ch0_timer_rst_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                       // CH0_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> CH0_TIMER_RST_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          ch0_timer_rst_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;               // CH0_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> CH0_TIMER_RST_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] ch0_timer_rst_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                        // CH0_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> CH0_TIMER_RST_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          ch0_timer_rst_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                       // CH0_TIMER_RST_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> CH0_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          ch0_timer_rst_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;              // CH0_TIMER_RST_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> CH0_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          ch0_timer_rst_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                    // CH0_TIMER_RST_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> CH0_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          ch0_timer_rst_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;            // CH0_TIMER_RST_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> CH0_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] ch0_timer_rst_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                     // CH0_TIMER_RST_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> CH0_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          ch0_timer_rst_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                    // CH0_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> CH0_TIMER_RST_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          ch0_timer_rst_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                  // CH0_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> CH0_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] ch0_timer_rst_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                   // CH0_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> CH0_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          ch0_timer_rst_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                  // CH0_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> CH0_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          detector_on_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                          // DETECTOR_ON_s1_translator:uav_waitrequest -> DETECTOR_ON_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] detector_on_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                           // DETECTOR_ON_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> DETECTOR_ON_s1_translator:uav_burstcount
	wire   [31:0] detector_on_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                            // DETECTOR_ON_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> DETECTOR_ON_s1_translator:uav_writedata
	wire   [21:0] detector_on_s1_translator_avalon_universal_slave_0_agent_m0_address;                              // DETECTOR_ON_s1_translator_avalon_universal_slave_0_agent:m0_address -> DETECTOR_ON_s1_translator:uav_address
	wire          detector_on_s1_translator_avalon_universal_slave_0_agent_m0_write;                                // DETECTOR_ON_s1_translator_avalon_universal_slave_0_agent:m0_write -> DETECTOR_ON_s1_translator:uav_write
	wire          detector_on_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                 // DETECTOR_ON_s1_translator_avalon_universal_slave_0_agent:m0_lock -> DETECTOR_ON_s1_translator:uav_lock
	wire          detector_on_s1_translator_avalon_universal_slave_0_agent_m0_read;                                 // DETECTOR_ON_s1_translator_avalon_universal_slave_0_agent:m0_read -> DETECTOR_ON_s1_translator:uav_read
	wire   [31:0] detector_on_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                             // DETECTOR_ON_s1_translator:uav_readdata -> DETECTOR_ON_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          detector_on_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                        // DETECTOR_ON_s1_translator:uav_readdatavalid -> DETECTOR_ON_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          detector_on_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                          // DETECTOR_ON_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> DETECTOR_ON_s1_translator:uav_debugaccess
	wire    [3:0] detector_on_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                           // DETECTOR_ON_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> DETECTOR_ON_s1_translator:uav_byteenable
	wire          detector_on_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                   // DETECTOR_ON_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> DETECTOR_ON_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          detector_on_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                         // DETECTOR_ON_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> DETECTOR_ON_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          detector_on_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                 // DETECTOR_ON_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> DETECTOR_ON_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] detector_on_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                          // DETECTOR_ON_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> DETECTOR_ON_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          detector_on_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                         // DETECTOR_ON_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> DETECTOR_ON_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          detector_on_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                // DETECTOR_ON_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> DETECTOR_ON_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          detector_on_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                      // DETECTOR_ON_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> DETECTOR_ON_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          detector_on_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;              // DETECTOR_ON_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> DETECTOR_ON_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] detector_on_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                       // DETECTOR_ON_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> DETECTOR_ON_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          detector_on_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                      // DETECTOR_ON_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> DETECTOR_ON_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          detector_on_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                    // DETECTOR_ON_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> DETECTOR_ON_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] detector_on_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                     // DETECTOR_ON_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> DETECTOR_ON_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          detector_on_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                    // DETECTOR_ON_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> DETECTOR_ON_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          menu_down_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                            // MENU_DOWN_s1_translator:uav_waitrequest -> MENU_DOWN_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] menu_down_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                             // MENU_DOWN_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> MENU_DOWN_s1_translator:uav_burstcount
	wire   [31:0] menu_down_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                              // MENU_DOWN_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> MENU_DOWN_s1_translator:uav_writedata
	wire   [21:0] menu_down_s1_translator_avalon_universal_slave_0_agent_m0_address;                                // MENU_DOWN_s1_translator_avalon_universal_slave_0_agent:m0_address -> MENU_DOWN_s1_translator:uav_address
	wire          menu_down_s1_translator_avalon_universal_slave_0_agent_m0_write;                                  // MENU_DOWN_s1_translator_avalon_universal_slave_0_agent:m0_write -> MENU_DOWN_s1_translator:uav_write
	wire          menu_down_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                   // MENU_DOWN_s1_translator_avalon_universal_slave_0_agent:m0_lock -> MENU_DOWN_s1_translator:uav_lock
	wire          menu_down_s1_translator_avalon_universal_slave_0_agent_m0_read;                                   // MENU_DOWN_s1_translator_avalon_universal_slave_0_agent:m0_read -> MENU_DOWN_s1_translator:uav_read
	wire   [31:0] menu_down_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                               // MENU_DOWN_s1_translator:uav_readdata -> MENU_DOWN_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          menu_down_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                          // MENU_DOWN_s1_translator:uav_readdatavalid -> MENU_DOWN_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          menu_down_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                            // MENU_DOWN_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> MENU_DOWN_s1_translator:uav_debugaccess
	wire    [3:0] menu_down_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                             // MENU_DOWN_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> MENU_DOWN_s1_translator:uav_byteenable
	wire          menu_down_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                     // MENU_DOWN_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> MENU_DOWN_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          menu_down_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                           // MENU_DOWN_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> MENU_DOWN_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          menu_down_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                   // MENU_DOWN_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> MENU_DOWN_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] menu_down_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                            // MENU_DOWN_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> MENU_DOWN_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          menu_down_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                           // MENU_DOWN_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> MENU_DOWN_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          menu_down_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                  // MENU_DOWN_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> MENU_DOWN_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          menu_down_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                        // MENU_DOWN_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> MENU_DOWN_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          menu_down_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                // MENU_DOWN_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> MENU_DOWN_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] menu_down_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                         // MENU_DOWN_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> MENU_DOWN_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          menu_down_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                        // MENU_DOWN_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> MENU_DOWN_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          menu_down_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                      // MENU_DOWN_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> MENU_DOWN_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] menu_down_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                       // MENU_DOWN_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> MENU_DOWN_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          menu_down_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                      // MENU_DOWN_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> MENU_DOWN_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          menu_up_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                              // MENU_UP_s1_translator:uav_waitrequest -> MENU_UP_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] menu_up_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                               // MENU_UP_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> MENU_UP_s1_translator:uav_burstcount
	wire   [31:0] menu_up_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                // MENU_UP_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> MENU_UP_s1_translator:uav_writedata
	wire   [21:0] menu_up_s1_translator_avalon_universal_slave_0_agent_m0_address;                                  // MENU_UP_s1_translator_avalon_universal_slave_0_agent:m0_address -> MENU_UP_s1_translator:uav_address
	wire          menu_up_s1_translator_avalon_universal_slave_0_agent_m0_write;                                    // MENU_UP_s1_translator_avalon_universal_slave_0_agent:m0_write -> MENU_UP_s1_translator:uav_write
	wire          menu_up_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                     // MENU_UP_s1_translator_avalon_universal_slave_0_agent:m0_lock -> MENU_UP_s1_translator:uav_lock
	wire          menu_up_s1_translator_avalon_universal_slave_0_agent_m0_read;                                     // MENU_UP_s1_translator_avalon_universal_slave_0_agent:m0_read -> MENU_UP_s1_translator:uav_read
	wire   [31:0] menu_up_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                 // MENU_UP_s1_translator:uav_readdata -> MENU_UP_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          menu_up_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                            // MENU_UP_s1_translator:uav_readdatavalid -> MENU_UP_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          menu_up_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                              // MENU_UP_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> MENU_UP_s1_translator:uav_debugaccess
	wire    [3:0] menu_up_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                               // MENU_UP_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> MENU_UP_s1_translator:uav_byteenable
	wire          menu_up_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                       // MENU_UP_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> MENU_UP_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          menu_up_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                             // MENU_UP_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> MENU_UP_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          menu_up_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                     // MENU_UP_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> MENU_UP_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] menu_up_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                              // MENU_UP_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> MENU_UP_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          menu_up_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                             // MENU_UP_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> MENU_UP_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          menu_up_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                    // MENU_UP_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> MENU_UP_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          menu_up_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                          // MENU_UP_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> MENU_UP_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          menu_up_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                  // MENU_UP_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> MENU_UP_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] menu_up_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                           // MENU_UP_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> MENU_UP_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          menu_up_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                          // MENU_UP_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> MENU_UP_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          menu_up_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                        // MENU_UP_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> MENU_UP_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] menu_up_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                         // MENU_UP_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> MENU_UP_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          menu_up_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                        // MENU_UP_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> MENU_UP_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          menu_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                 // MENU_s1_translator:uav_waitrequest -> MENU_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] menu_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                  // MENU_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> MENU_s1_translator:uav_burstcount
	wire   [31:0] menu_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                   // MENU_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> MENU_s1_translator:uav_writedata
	wire   [21:0] menu_s1_translator_avalon_universal_slave_0_agent_m0_address;                                     // MENU_s1_translator_avalon_universal_slave_0_agent:m0_address -> MENU_s1_translator:uav_address
	wire          menu_s1_translator_avalon_universal_slave_0_agent_m0_write;                                       // MENU_s1_translator_avalon_universal_slave_0_agent:m0_write -> MENU_s1_translator:uav_write
	wire          menu_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                        // MENU_s1_translator_avalon_universal_slave_0_agent:m0_lock -> MENU_s1_translator:uav_lock
	wire          menu_s1_translator_avalon_universal_slave_0_agent_m0_read;                                        // MENU_s1_translator_avalon_universal_slave_0_agent:m0_read -> MENU_s1_translator:uav_read
	wire   [31:0] menu_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                    // MENU_s1_translator:uav_readdata -> MENU_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          menu_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                               // MENU_s1_translator:uav_readdatavalid -> MENU_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          menu_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                 // MENU_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> MENU_s1_translator:uav_debugaccess
	wire    [3:0] menu_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                  // MENU_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> MENU_s1_translator:uav_byteenable
	wire          menu_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                          // MENU_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> MENU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          menu_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                // MENU_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> MENU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          menu_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                        // MENU_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> MENU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] menu_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                 // MENU_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> MENU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          menu_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                // MENU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> MENU_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          menu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                       // MENU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> MENU_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          menu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                             // MENU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> MENU_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          menu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                     // MENU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> MENU_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] menu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                              // MENU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> MENU_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          menu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                             // MENU_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> MENU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          menu_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                           // MENU_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> MENU_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] menu_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                            // MENU_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> MENU_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          menu_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                           // MENU_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> MENU_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          ch0_thresh_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                           // CH0_THRESH_s1_translator:uav_waitrequest -> CH0_THRESH_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] ch0_thresh_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                            // CH0_THRESH_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> CH0_THRESH_s1_translator:uav_burstcount
	wire   [31:0] ch0_thresh_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                             // CH0_THRESH_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> CH0_THRESH_s1_translator:uav_writedata
	wire   [21:0] ch0_thresh_s1_translator_avalon_universal_slave_0_agent_m0_address;                               // CH0_THRESH_s1_translator_avalon_universal_slave_0_agent:m0_address -> CH0_THRESH_s1_translator:uav_address
	wire          ch0_thresh_s1_translator_avalon_universal_slave_0_agent_m0_write;                                 // CH0_THRESH_s1_translator_avalon_universal_slave_0_agent:m0_write -> CH0_THRESH_s1_translator:uav_write
	wire          ch0_thresh_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                  // CH0_THRESH_s1_translator_avalon_universal_slave_0_agent:m0_lock -> CH0_THRESH_s1_translator:uav_lock
	wire          ch0_thresh_s1_translator_avalon_universal_slave_0_agent_m0_read;                                  // CH0_THRESH_s1_translator_avalon_universal_slave_0_agent:m0_read -> CH0_THRESH_s1_translator:uav_read
	wire   [31:0] ch0_thresh_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                              // CH0_THRESH_s1_translator:uav_readdata -> CH0_THRESH_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          ch0_thresh_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                         // CH0_THRESH_s1_translator:uav_readdatavalid -> CH0_THRESH_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          ch0_thresh_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                           // CH0_THRESH_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> CH0_THRESH_s1_translator:uav_debugaccess
	wire    [3:0] ch0_thresh_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                            // CH0_THRESH_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> CH0_THRESH_s1_translator:uav_byteenable
	wire          ch0_thresh_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                    // CH0_THRESH_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> CH0_THRESH_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          ch0_thresh_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                          // CH0_THRESH_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> CH0_THRESH_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          ch0_thresh_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                  // CH0_THRESH_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> CH0_THRESH_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] ch0_thresh_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                           // CH0_THRESH_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> CH0_THRESH_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          ch0_thresh_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                          // CH0_THRESH_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> CH0_THRESH_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          ch0_thresh_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                 // CH0_THRESH_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> CH0_THRESH_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          ch0_thresh_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                       // CH0_THRESH_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> CH0_THRESH_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          ch0_thresh_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;               // CH0_THRESH_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> CH0_THRESH_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] ch0_thresh_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                        // CH0_THRESH_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> CH0_THRESH_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          ch0_thresh_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                       // CH0_THRESH_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> CH0_THRESH_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          ch0_thresh_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                     // CH0_THRESH_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> CH0_THRESH_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] ch0_thresh_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                      // CH0_THRESH_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> CH0_THRESH_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          ch0_thresh_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                     // CH0_THRESH_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> CH0_THRESH_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          ch0_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                          // CH0_RD_PEAK_s1_translator:uav_waitrequest -> CH0_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] ch0_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                           // CH0_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> CH0_RD_PEAK_s1_translator:uav_burstcount
	wire   [31:0] ch0_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                            // CH0_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> CH0_RD_PEAK_s1_translator:uav_writedata
	wire   [21:0] ch0_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_address;                              // CH0_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:m0_address -> CH0_RD_PEAK_s1_translator:uav_address
	wire          ch0_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_write;                                // CH0_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:m0_write -> CH0_RD_PEAK_s1_translator:uav_write
	wire          ch0_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                 // CH0_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:m0_lock -> CH0_RD_PEAK_s1_translator:uav_lock
	wire          ch0_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_read;                                 // CH0_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:m0_read -> CH0_RD_PEAK_s1_translator:uav_read
	wire   [31:0] ch0_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                             // CH0_RD_PEAK_s1_translator:uav_readdata -> CH0_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          ch0_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                        // CH0_RD_PEAK_s1_translator:uav_readdatavalid -> CH0_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          ch0_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                          // CH0_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> CH0_RD_PEAK_s1_translator:uav_debugaccess
	wire    [3:0] ch0_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                           // CH0_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> CH0_RD_PEAK_s1_translator:uav_byteenable
	wire          ch0_rd_peak_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                   // CH0_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> CH0_RD_PEAK_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          ch0_rd_peak_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                         // CH0_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> CH0_RD_PEAK_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          ch0_rd_peak_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                 // CH0_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> CH0_RD_PEAK_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] ch0_rd_peak_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                          // CH0_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> CH0_RD_PEAK_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          ch0_rd_peak_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                         // CH0_RD_PEAK_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> CH0_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          ch0_rd_peak_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                // CH0_RD_PEAK_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> CH0_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          ch0_rd_peak_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                      // CH0_RD_PEAK_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> CH0_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          ch0_rd_peak_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;              // CH0_RD_PEAK_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> CH0_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] ch0_rd_peak_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                       // CH0_RD_PEAK_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> CH0_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          ch0_rd_peak_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                      // CH0_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> CH0_RD_PEAK_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          ch0_rd_peak_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                    // CH0_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> CH0_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] ch0_rd_peak_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                     // CH0_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> CH0_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          ch0_rd_peak_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                    // CH0_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> CH0_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          ch0_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                       // CH0_PEAK_FOUND_s1_translator:uav_waitrequest -> CH0_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] ch0_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                        // CH0_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> CH0_PEAK_FOUND_s1_translator:uav_burstcount
	wire   [31:0] ch0_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                         // CH0_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> CH0_PEAK_FOUND_s1_translator:uav_writedata
	wire   [21:0] ch0_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_address;                           // CH0_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:m0_address -> CH0_PEAK_FOUND_s1_translator:uav_address
	wire          ch0_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_write;                             // CH0_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:m0_write -> CH0_PEAK_FOUND_s1_translator:uav_write
	wire          ch0_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_lock;                              // CH0_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:m0_lock -> CH0_PEAK_FOUND_s1_translator:uav_lock
	wire          ch0_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_read;                              // CH0_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:m0_read -> CH0_PEAK_FOUND_s1_translator:uav_read
	wire   [31:0] ch0_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                          // CH0_PEAK_FOUND_s1_translator:uav_readdata -> CH0_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          ch0_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                     // CH0_PEAK_FOUND_s1_translator:uav_readdatavalid -> CH0_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          ch0_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                       // CH0_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> CH0_PEAK_FOUND_s1_translator:uav_debugaccess
	wire    [3:0] ch0_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                        // CH0_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> CH0_PEAK_FOUND_s1_translator:uav_byteenable
	wire          ch0_peak_found_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                // CH0_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> CH0_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          ch0_peak_found_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                      // CH0_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> CH0_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          ch0_peak_found_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;              // CH0_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> CH0_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] ch0_peak_found_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                       // CH0_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> CH0_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          ch0_peak_found_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                      // CH0_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> CH0_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          ch0_peak_found_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;             // CH0_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> CH0_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          ch0_peak_found_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                   // CH0_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> CH0_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          ch0_peak_found_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;           // CH0_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> CH0_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] ch0_peak_found_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                    // CH0_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> CH0_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          ch0_peak_found_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                   // CH0_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> CH0_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          ch0_peak_found_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                 // CH0_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> CH0_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] ch0_peak_found_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                  // CH0_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> CH0_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          ch0_peak_found_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                 // CH0_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> CH0_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          ch0_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                            // CH0_YN1_L_s1_translator:uav_waitrequest -> CH0_YN1_L_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] ch0_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                             // CH0_YN1_L_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> CH0_YN1_L_s1_translator:uav_burstcount
	wire   [31:0] ch0_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                              // CH0_YN1_L_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> CH0_YN1_L_s1_translator:uav_writedata
	wire   [21:0] ch0_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_address;                                // CH0_YN1_L_s1_translator_avalon_universal_slave_0_agent:m0_address -> CH0_YN1_L_s1_translator:uav_address
	wire          ch0_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_write;                                  // CH0_YN1_L_s1_translator_avalon_universal_slave_0_agent:m0_write -> CH0_YN1_L_s1_translator:uav_write
	wire          ch0_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                   // CH0_YN1_L_s1_translator_avalon_universal_slave_0_agent:m0_lock -> CH0_YN1_L_s1_translator:uav_lock
	wire          ch0_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_read;                                   // CH0_YN1_L_s1_translator_avalon_universal_slave_0_agent:m0_read -> CH0_YN1_L_s1_translator:uav_read
	wire   [31:0] ch0_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                               // CH0_YN1_L_s1_translator:uav_readdata -> CH0_YN1_L_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          ch0_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                          // CH0_YN1_L_s1_translator:uav_readdatavalid -> CH0_YN1_L_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          ch0_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                            // CH0_YN1_L_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> CH0_YN1_L_s1_translator:uav_debugaccess
	wire    [3:0] ch0_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                             // CH0_YN1_L_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> CH0_YN1_L_s1_translator:uav_byteenable
	wire          ch0_yn1_l_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                     // CH0_YN1_L_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> CH0_YN1_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          ch0_yn1_l_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                           // CH0_YN1_L_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> CH0_YN1_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          ch0_yn1_l_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                   // CH0_YN1_L_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> CH0_YN1_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] ch0_yn1_l_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                            // CH0_YN1_L_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> CH0_YN1_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          ch0_yn1_l_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                           // CH0_YN1_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> CH0_YN1_L_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          ch0_yn1_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                  // CH0_YN1_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> CH0_YN1_L_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          ch0_yn1_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                        // CH0_YN1_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> CH0_YN1_L_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          ch0_yn1_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                // CH0_YN1_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> CH0_YN1_L_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] ch0_yn1_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                         // CH0_YN1_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> CH0_YN1_L_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          ch0_yn1_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                        // CH0_YN1_L_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> CH0_YN1_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          ch0_yn1_l_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                      // CH0_YN1_L_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> CH0_YN1_L_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] ch0_yn1_l_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                       // CH0_YN1_L_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> CH0_YN1_L_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          ch0_yn1_l_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                      // CH0_YN1_L_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> CH0_YN1_L_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          ch0_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                           // CH0_YN1_ML_s1_translator:uav_waitrequest -> CH0_YN1_ML_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] ch0_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                            // CH0_YN1_ML_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> CH0_YN1_ML_s1_translator:uav_burstcount
	wire   [31:0] ch0_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                             // CH0_YN1_ML_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> CH0_YN1_ML_s1_translator:uav_writedata
	wire   [21:0] ch0_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_address;                               // CH0_YN1_ML_s1_translator_avalon_universal_slave_0_agent:m0_address -> CH0_YN1_ML_s1_translator:uav_address
	wire          ch0_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_write;                                 // CH0_YN1_ML_s1_translator_avalon_universal_slave_0_agent:m0_write -> CH0_YN1_ML_s1_translator:uav_write
	wire          ch0_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                  // CH0_YN1_ML_s1_translator_avalon_universal_slave_0_agent:m0_lock -> CH0_YN1_ML_s1_translator:uav_lock
	wire          ch0_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_read;                                  // CH0_YN1_ML_s1_translator_avalon_universal_slave_0_agent:m0_read -> CH0_YN1_ML_s1_translator:uav_read
	wire   [31:0] ch0_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                              // CH0_YN1_ML_s1_translator:uav_readdata -> CH0_YN1_ML_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          ch0_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                         // CH0_YN1_ML_s1_translator:uav_readdatavalid -> CH0_YN1_ML_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          ch0_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                           // CH0_YN1_ML_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> CH0_YN1_ML_s1_translator:uav_debugaccess
	wire    [3:0] ch0_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                            // CH0_YN1_ML_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> CH0_YN1_ML_s1_translator:uav_byteenable
	wire          ch0_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                    // CH0_YN1_ML_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> CH0_YN1_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          ch0_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                          // CH0_YN1_ML_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> CH0_YN1_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          ch0_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                  // CH0_YN1_ML_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> CH0_YN1_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] ch0_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                           // CH0_YN1_ML_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> CH0_YN1_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          ch0_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                          // CH0_YN1_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> CH0_YN1_ML_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          ch0_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                 // CH0_YN1_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> CH0_YN1_ML_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          ch0_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                       // CH0_YN1_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> CH0_YN1_ML_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          ch0_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;               // CH0_YN1_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> CH0_YN1_ML_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] ch0_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                        // CH0_YN1_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> CH0_YN1_ML_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          ch0_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                       // CH0_YN1_ML_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> CH0_YN1_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          ch0_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                     // CH0_YN1_ML_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> CH0_YN1_ML_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] ch0_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                      // CH0_YN1_ML_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> CH0_YN1_ML_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          ch0_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                     // CH0_YN1_ML_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> CH0_YN1_ML_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          ch0_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                           // CH0_YN1_MU_s1_translator:uav_waitrequest -> CH0_YN1_MU_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] ch0_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                            // CH0_YN1_MU_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> CH0_YN1_MU_s1_translator:uav_burstcount
	wire   [31:0] ch0_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                             // CH0_YN1_MU_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> CH0_YN1_MU_s1_translator:uav_writedata
	wire   [21:0] ch0_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_address;                               // CH0_YN1_MU_s1_translator_avalon_universal_slave_0_agent:m0_address -> CH0_YN1_MU_s1_translator:uav_address
	wire          ch0_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_write;                                 // CH0_YN1_MU_s1_translator_avalon_universal_slave_0_agent:m0_write -> CH0_YN1_MU_s1_translator:uav_write
	wire          ch0_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                  // CH0_YN1_MU_s1_translator_avalon_universal_slave_0_agent:m0_lock -> CH0_YN1_MU_s1_translator:uav_lock
	wire          ch0_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_read;                                  // CH0_YN1_MU_s1_translator_avalon_universal_slave_0_agent:m0_read -> CH0_YN1_MU_s1_translator:uav_read
	wire   [31:0] ch0_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                              // CH0_YN1_MU_s1_translator:uav_readdata -> CH0_YN1_MU_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          ch0_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                         // CH0_YN1_MU_s1_translator:uav_readdatavalid -> CH0_YN1_MU_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          ch0_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                           // CH0_YN1_MU_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> CH0_YN1_MU_s1_translator:uav_debugaccess
	wire    [3:0] ch0_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                            // CH0_YN1_MU_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> CH0_YN1_MU_s1_translator:uav_byteenable
	wire          ch0_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                    // CH0_YN1_MU_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> CH0_YN1_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          ch0_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                          // CH0_YN1_MU_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> CH0_YN1_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          ch0_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                  // CH0_YN1_MU_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> CH0_YN1_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] ch0_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                           // CH0_YN1_MU_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> CH0_YN1_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          ch0_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                          // CH0_YN1_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> CH0_YN1_MU_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          ch0_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                 // CH0_YN1_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> CH0_YN1_MU_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          ch0_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                       // CH0_YN1_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> CH0_YN1_MU_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          ch0_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;               // CH0_YN1_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> CH0_YN1_MU_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] ch0_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                        // CH0_YN1_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> CH0_YN1_MU_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          ch0_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                       // CH0_YN1_MU_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> CH0_YN1_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          ch0_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                     // CH0_YN1_MU_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> CH0_YN1_MU_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] ch0_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                      // CH0_YN1_MU_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> CH0_YN1_MU_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          ch0_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                     // CH0_YN1_MU_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> CH0_YN1_MU_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          ch0_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                            // CH0_YN1_U_s1_translator:uav_waitrequest -> CH0_YN1_U_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] ch0_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                             // CH0_YN1_U_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> CH0_YN1_U_s1_translator:uav_burstcount
	wire   [31:0] ch0_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                              // CH0_YN1_U_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> CH0_YN1_U_s1_translator:uav_writedata
	wire   [21:0] ch0_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_address;                                // CH0_YN1_U_s1_translator_avalon_universal_slave_0_agent:m0_address -> CH0_YN1_U_s1_translator:uav_address
	wire          ch0_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_write;                                  // CH0_YN1_U_s1_translator_avalon_universal_slave_0_agent:m0_write -> CH0_YN1_U_s1_translator:uav_write
	wire          ch0_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                   // CH0_YN1_U_s1_translator_avalon_universal_slave_0_agent:m0_lock -> CH0_YN1_U_s1_translator:uav_lock
	wire          ch0_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_read;                                   // CH0_YN1_U_s1_translator_avalon_universal_slave_0_agent:m0_read -> CH0_YN1_U_s1_translator:uav_read
	wire   [31:0] ch0_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                               // CH0_YN1_U_s1_translator:uav_readdata -> CH0_YN1_U_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          ch0_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                          // CH0_YN1_U_s1_translator:uav_readdatavalid -> CH0_YN1_U_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          ch0_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                            // CH0_YN1_U_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> CH0_YN1_U_s1_translator:uav_debugaccess
	wire    [3:0] ch0_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                             // CH0_YN1_U_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> CH0_YN1_U_s1_translator:uav_byteenable
	wire          ch0_yn1_u_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                     // CH0_YN1_U_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> CH0_YN1_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          ch0_yn1_u_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                           // CH0_YN1_U_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> CH0_YN1_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          ch0_yn1_u_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                   // CH0_YN1_U_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> CH0_YN1_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] ch0_yn1_u_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                            // CH0_YN1_U_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> CH0_YN1_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          ch0_yn1_u_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                           // CH0_YN1_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> CH0_YN1_U_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          ch0_yn1_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                  // CH0_YN1_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> CH0_YN1_U_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          ch0_yn1_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                        // CH0_YN1_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> CH0_YN1_U_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          ch0_yn1_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                // CH0_YN1_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> CH0_YN1_U_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] ch0_yn1_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                         // CH0_YN1_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> CH0_YN1_U_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          ch0_yn1_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                        // CH0_YN1_U_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> CH0_YN1_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          ch0_yn1_u_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                      // CH0_YN1_U_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> CH0_YN1_U_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] ch0_yn1_u_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                       // CH0_YN1_U_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> CH0_YN1_U_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          ch0_yn1_u_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                      // CH0_YN1_U_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> CH0_YN1_U_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          ch0_time_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                             // CH0_TIME_s1_translator:uav_waitrequest -> CH0_TIME_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] ch0_time_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                              // CH0_TIME_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> CH0_TIME_s1_translator:uav_burstcount
	wire   [31:0] ch0_time_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                               // CH0_TIME_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> CH0_TIME_s1_translator:uav_writedata
	wire   [21:0] ch0_time_s1_translator_avalon_universal_slave_0_agent_m0_address;                                 // CH0_TIME_s1_translator_avalon_universal_slave_0_agent:m0_address -> CH0_TIME_s1_translator:uav_address
	wire          ch0_time_s1_translator_avalon_universal_slave_0_agent_m0_write;                                   // CH0_TIME_s1_translator_avalon_universal_slave_0_agent:m0_write -> CH0_TIME_s1_translator:uav_write
	wire          ch0_time_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                    // CH0_TIME_s1_translator_avalon_universal_slave_0_agent:m0_lock -> CH0_TIME_s1_translator:uav_lock
	wire          ch0_time_s1_translator_avalon_universal_slave_0_agent_m0_read;                                    // CH0_TIME_s1_translator_avalon_universal_slave_0_agent:m0_read -> CH0_TIME_s1_translator:uav_read
	wire   [31:0] ch0_time_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                // CH0_TIME_s1_translator:uav_readdata -> CH0_TIME_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          ch0_time_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                           // CH0_TIME_s1_translator:uav_readdatavalid -> CH0_TIME_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          ch0_time_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                             // CH0_TIME_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> CH0_TIME_s1_translator:uav_debugaccess
	wire    [3:0] ch0_time_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                              // CH0_TIME_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> CH0_TIME_s1_translator:uav_byteenable
	wire          ch0_time_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                      // CH0_TIME_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> CH0_TIME_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          ch0_time_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                            // CH0_TIME_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> CH0_TIME_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          ch0_time_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                    // CH0_TIME_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> CH0_TIME_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] ch0_time_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                             // CH0_TIME_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> CH0_TIME_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          ch0_time_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                            // CH0_TIME_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> CH0_TIME_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          ch0_time_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                   // CH0_TIME_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> CH0_TIME_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          ch0_time_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                         // CH0_TIME_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> CH0_TIME_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          ch0_time_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                 // CH0_TIME_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> CH0_TIME_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] ch0_time_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                          // CH0_TIME_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> CH0_TIME_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          ch0_time_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                         // CH0_TIME_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> CH0_TIME_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          ch0_time_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                       // CH0_TIME_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> CH0_TIME_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] ch0_time_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                        // CH0_TIME_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> CH0_TIME_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          ch0_time_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                       // CH0_TIME_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> CH0_TIME_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          ch0_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                           // CH0_YN2_MU_s1_translator:uav_waitrequest -> CH0_YN2_MU_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] ch0_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                            // CH0_YN2_MU_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> CH0_YN2_MU_s1_translator:uav_burstcount
	wire   [31:0] ch0_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                             // CH0_YN2_MU_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> CH0_YN2_MU_s1_translator:uav_writedata
	wire   [21:0] ch0_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_address;                               // CH0_YN2_MU_s1_translator_avalon_universal_slave_0_agent:m0_address -> CH0_YN2_MU_s1_translator:uav_address
	wire          ch0_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_write;                                 // CH0_YN2_MU_s1_translator_avalon_universal_slave_0_agent:m0_write -> CH0_YN2_MU_s1_translator:uav_write
	wire          ch0_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                  // CH0_YN2_MU_s1_translator_avalon_universal_slave_0_agent:m0_lock -> CH0_YN2_MU_s1_translator:uav_lock
	wire          ch0_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_read;                                  // CH0_YN2_MU_s1_translator_avalon_universal_slave_0_agent:m0_read -> CH0_YN2_MU_s1_translator:uav_read
	wire   [31:0] ch0_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                              // CH0_YN2_MU_s1_translator:uav_readdata -> CH0_YN2_MU_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          ch0_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                         // CH0_YN2_MU_s1_translator:uav_readdatavalid -> CH0_YN2_MU_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          ch0_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                           // CH0_YN2_MU_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> CH0_YN2_MU_s1_translator:uav_debugaccess
	wire    [3:0] ch0_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                            // CH0_YN2_MU_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> CH0_YN2_MU_s1_translator:uav_byteenable
	wire          ch0_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                    // CH0_YN2_MU_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> CH0_YN2_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          ch0_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                          // CH0_YN2_MU_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> CH0_YN2_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          ch0_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                  // CH0_YN2_MU_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> CH0_YN2_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] ch0_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                           // CH0_YN2_MU_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> CH0_YN2_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          ch0_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                          // CH0_YN2_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> CH0_YN2_MU_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          ch0_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                 // CH0_YN2_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> CH0_YN2_MU_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          ch0_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                       // CH0_YN2_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> CH0_YN2_MU_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          ch0_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;               // CH0_YN2_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> CH0_YN2_MU_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] ch0_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                        // CH0_YN2_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> CH0_YN2_MU_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          ch0_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                       // CH0_YN2_MU_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> CH0_YN2_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          ch0_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                     // CH0_YN2_MU_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> CH0_YN2_MU_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] ch0_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                      // CH0_YN2_MU_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> CH0_YN2_MU_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          ch0_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                     // CH0_YN2_MU_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> CH0_YN2_MU_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          ch0_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                           // CH0_YN2_ML_s1_translator:uav_waitrequest -> CH0_YN2_ML_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] ch0_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                            // CH0_YN2_ML_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> CH0_YN2_ML_s1_translator:uav_burstcount
	wire   [31:0] ch0_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                             // CH0_YN2_ML_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> CH0_YN2_ML_s1_translator:uav_writedata
	wire   [21:0] ch0_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_address;                               // CH0_YN2_ML_s1_translator_avalon_universal_slave_0_agent:m0_address -> CH0_YN2_ML_s1_translator:uav_address
	wire          ch0_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_write;                                 // CH0_YN2_ML_s1_translator_avalon_universal_slave_0_agent:m0_write -> CH0_YN2_ML_s1_translator:uav_write
	wire          ch0_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                  // CH0_YN2_ML_s1_translator_avalon_universal_slave_0_agent:m0_lock -> CH0_YN2_ML_s1_translator:uav_lock
	wire          ch0_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_read;                                  // CH0_YN2_ML_s1_translator_avalon_universal_slave_0_agent:m0_read -> CH0_YN2_ML_s1_translator:uav_read
	wire   [31:0] ch0_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                              // CH0_YN2_ML_s1_translator:uav_readdata -> CH0_YN2_ML_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          ch0_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                         // CH0_YN2_ML_s1_translator:uav_readdatavalid -> CH0_YN2_ML_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          ch0_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                           // CH0_YN2_ML_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> CH0_YN2_ML_s1_translator:uav_debugaccess
	wire    [3:0] ch0_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                            // CH0_YN2_ML_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> CH0_YN2_ML_s1_translator:uav_byteenable
	wire          ch0_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                    // CH0_YN2_ML_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> CH0_YN2_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          ch0_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                          // CH0_YN2_ML_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> CH0_YN2_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          ch0_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                  // CH0_YN2_ML_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> CH0_YN2_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] ch0_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                           // CH0_YN2_ML_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> CH0_YN2_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          ch0_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                          // CH0_YN2_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> CH0_YN2_ML_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          ch0_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                 // CH0_YN2_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> CH0_YN2_ML_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          ch0_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                       // CH0_YN2_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> CH0_YN2_ML_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          ch0_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;               // CH0_YN2_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> CH0_YN2_ML_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] ch0_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                        // CH0_YN2_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> CH0_YN2_ML_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          ch0_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                       // CH0_YN2_ML_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> CH0_YN2_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          ch0_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                     // CH0_YN2_ML_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> CH0_YN2_ML_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] ch0_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                      // CH0_YN2_ML_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> CH0_YN2_ML_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          ch0_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                     // CH0_YN2_ML_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> CH0_YN2_ML_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          ch0_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                            // CH0_YN2_U_s1_translator:uav_waitrequest -> CH0_YN2_U_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] ch0_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                             // CH0_YN2_U_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> CH0_YN2_U_s1_translator:uav_burstcount
	wire   [31:0] ch0_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                              // CH0_YN2_U_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> CH0_YN2_U_s1_translator:uav_writedata
	wire   [21:0] ch0_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_address;                                // CH0_YN2_U_s1_translator_avalon_universal_slave_0_agent:m0_address -> CH0_YN2_U_s1_translator:uav_address
	wire          ch0_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_write;                                  // CH0_YN2_U_s1_translator_avalon_universal_slave_0_agent:m0_write -> CH0_YN2_U_s1_translator:uav_write
	wire          ch0_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                   // CH0_YN2_U_s1_translator_avalon_universal_slave_0_agent:m0_lock -> CH0_YN2_U_s1_translator:uav_lock
	wire          ch0_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_read;                                   // CH0_YN2_U_s1_translator_avalon_universal_slave_0_agent:m0_read -> CH0_YN2_U_s1_translator:uav_read
	wire   [31:0] ch0_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                               // CH0_YN2_U_s1_translator:uav_readdata -> CH0_YN2_U_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          ch0_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                          // CH0_YN2_U_s1_translator:uav_readdatavalid -> CH0_YN2_U_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          ch0_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                            // CH0_YN2_U_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> CH0_YN2_U_s1_translator:uav_debugaccess
	wire    [3:0] ch0_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                             // CH0_YN2_U_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> CH0_YN2_U_s1_translator:uav_byteenable
	wire          ch0_yn2_u_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                     // CH0_YN2_U_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> CH0_YN2_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          ch0_yn2_u_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                           // CH0_YN2_U_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> CH0_YN2_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          ch0_yn2_u_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                   // CH0_YN2_U_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> CH0_YN2_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] ch0_yn2_u_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                            // CH0_YN2_U_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> CH0_YN2_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          ch0_yn2_u_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                           // CH0_YN2_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> CH0_YN2_U_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          ch0_yn2_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                  // CH0_YN2_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> CH0_YN2_U_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          ch0_yn2_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                        // CH0_YN2_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> CH0_YN2_U_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          ch0_yn2_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                // CH0_YN2_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> CH0_YN2_U_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] ch0_yn2_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                         // CH0_YN2_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> CH0_YN2_U_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          ch0_yn2_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                        // CH0_YN2_U_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> CH0_YN2_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          ch0_yn2_u_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                      // CH0_YN2_U_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> CH0_YN2_U_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] ch0_yn2_u_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                       // CH0_YN2_U_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> CH0_YN2_U_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          ch0_yn2_u_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                      // CH0_YN2_U_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> CH0_YN2_U_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          ch0_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                            // CH0_YN2_L_s1_translator:uav_waitrequest -> CH0_YN2_L_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] ch0_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                             // CH0_YN2_L_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> CH0_YN2_L_s1_translator:uav_burstcount
	wire   [31:0] ch0_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                              // CH0_YN2_L_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> CH0_YN2_L_s1_translator:uav_writedata
	wire   [21:0] ch0_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_address;                                // CH0_YN2_L_s1_translator_avalon_universal_slave_0_agent:m0_address -> CH0_YN2_L_s1_translator:uav_address
	wire          ch0_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_write;                                  // CH0_YN2_L_s1_translator_avalon_universal_slave_0_agent:m0_write -> CH0_YN2_L_s1_translator:uav_write
	wire          ch0_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                   // CH0_YN2_L_s1_translator_avalon_universal_slave_0_agent:m0_lock -> CH0_YN2_L_s1_translator:uav_lock
	wire          ch0_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_read;                                   // CH0_YN2_L_s1_translator_avalon_universal_slave_0_agent:m0_read -> CH0_YN2_L_s1_translator:uav_read
	wire   [31:0] ch0_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                               // CH0_YN2_L_s1_translator:uav_readdata -> CH0_YN2_L_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          ch0_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                          // CH0_YN2_L_s1_translator:uav_readdatavalid -> CH0_YN2_L_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          ch0_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                            // CH0_YN2_L_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> CH0_YN2_L_s1_translator:uav_debugaccess
	wire    [3:0] ch0_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                             // CH0_YN2_L_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> CH0_YN2_L_s1_translator:uav_byteenable
	wire          ch0_yn2_l_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                     // CH0_YN2_L_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> CH0_YN2_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          ch0_yn2_l_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                           // CH0_YN2_L_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> CH0_YN2_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          ch0_yn2_l_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                   // CH0_YN2_L_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> CH0_YN2_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] ch0_yn2_l_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                            // CH0_YN2_L_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> CH0_YN2_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          ch0_yn2_l_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                           // CH0_YN2_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> CH0_YN2_L_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          ch0_yn2_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                  // CH0_YN2_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> CH0_YN2_L_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          ch0_yn2_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                        // CH0_YN2_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> CH0_YN2_L_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          ch0_yn2_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                // CH0_YN2_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> CH0_YN2_L_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] ch0_yn2_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                         // CH0_YN2_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> CH0_YN2_L_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          ch0_yn2_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                        // CH0_YN2_L_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> CH0_YN2_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          ch0_yn2_l_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                      // CH0_YN2_L_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> CH0_YN2_L_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] ch0_yn2_l_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                       // CH0_YN2_L_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> CH0_YN2_L_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          ch0_yn2_l_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                      // CH0_YN2_L_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> CH0_YN2_L_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          ch0_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                            // CH0_YN3_L_s1_translator:uav_waitrequest -> CH0_YN3_L_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] ch0_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                             // CH0_YN3_L_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> CH0_YN3_L_s1_translator:uav_burstcount
	wire   [31:0] ch0_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                              // CH0_YN3_L_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> CH0_YN3_L_s1_translator:uav_writedata
	wire   [21:0] ch0_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_address;                                // CH0_YN3_L_s1_translator_avalon_universal_slave_0_agent:m0_address -> CH0_YN3_L_s1_translator:uav_address
	wire          ch0_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_write;                                  // CH0_YN3_L_s1_translator_avalon_universal_slave_0_agent:m0_write -> CH0_YN3_L_s1_translator:uav_write
	wire          ch0_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                   // CH0_YN3_L_s1_translator_avalon_universal_slave_0_agent:m0_lock -> CH0_YN3_L_s1_translator:uav_lock
	wire          ch0_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_read;                                   // CH0_YN3_L_s1_translator_avalon_universal_slave_0_agent:m0_read -> CH0_YN3_L_s1_translator:uav_read
	wire   [31:0] ch0_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                               // CH0_YN3_L_s1_translator:uav_readdata -> CH0_YN3_L_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          ch0_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                          // CH0_YN3_L_s1_translator:uav_readdatavalid -> CH0_YN3_L_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          ch0_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                            // CH0_YN3_L_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> CH0_YN3_L_s1_translator:uav_debugaccess
	wire    [3:0] ch0_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                             // CH0_YN3_L_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> CH0_YN3_L_s1_translator:uav_byteenable
	wire          ch0_yn3_l_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                     // CH0_YN3_L_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> CH0_YN3_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          ch0_yn3_l_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                           // CH0_YN3_L_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> CH0_YN3_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          ch0_yn3_l_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                   // CH0_YN3_L_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> CH0_YN3_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] ch0_yn3_l_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                            // CH0_YN3_L_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> CH0_YN3_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          ch0_yn3_l_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                           // CH0_YN3_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> CH0_YN3_L_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          ch0_yn3_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                  // CH0_YN3_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> CH0_YN3_L_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          ch0_yn3_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                        // CH0_YN3_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> CH0_YN3_L_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          ch0_yn3_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                // CH0_YN3_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> CH0_YN3_L_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] ch0_yn3_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                         // CH0_YN3_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> CH0_YN3_L_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          ch0_yn3_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                        // CH0_YN3_L_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> CH0_YN3_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          ch0_yn3_l_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                      // CH0_YN3_L_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> CH0_YN3_L_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] ch0_yn3_l_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                       // CH0_YN3_L_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> CH0_YN3_L_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          ch0_yn3_l_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                      // CH0_YN3_L_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> CH0_YN3_L_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          ch0_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                           // CH0_YN3_ML_s1_translator:uav_waitrequest -> CH0_YN3_ML_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] ch0_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                            // CH0_YN3_ML_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> CH0_YN3_ML_s1_translator:uav_burstcount
	wire   [31:0] ch0_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                             // CH0_YN3_ML_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> CH0_YN3_ML_s1_translator:uav_writedata
	wire   [21:0] ch0_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_address;                               // CH0_YN3_ML_s1_translator_avalon_universal_slave_0_agent:m0_address -> CH0_YN3_ML_s1_translator:uav_address
	wire          ch0_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_write;                                 // CH0_YN3_ML_s1_translator_avalon_universal_slave_0_agent:m0_write -> CH0_YN3_ML_s1_translator:uav_write
	wire          ch0_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                  // CH0_YN3_ML_s1_translator_avalon_universal_slave_0_agent:m0_lock -> CH0_YN3_ML_s1_translator:uav_lock
	wire          ch0_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_read;                                  // CH0_YN3_ML_s1_translator_avalon_universal_slave_0_agent:m0_read -> CH0_YN3_ML_s1_translator:uav_read
	wire   [31:0] ch0_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                              // CH0_YN3_ML_s1_translator:uav_readdata -> CH0_YN3_ML_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          ch0_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                         // CH0_YN3_ML_s1_translator:uav_readdatavalid -> CH0_YN3_ML_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          ch0_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                           // CH0_YN3_ML_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> CH0_YN3_ML_s1_translator:uav_debugaccess
	wire    [3:0] ch0_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                            // CH0_YN3_ML_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> CH0_YN3_ML_s1_translator:uav_byteenable
	wire          ch0_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                    // CH0_YN3_ML_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> CH0_YN3_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          ch0_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                          // CH0_YN3_ML_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> CH0_YN3_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          ch0_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                  // CH0_YN3_ML_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> CH0_YN3_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] ch0_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                           // CH0_YN3_ML_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> CH0_YN3_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          ch0_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                          // CH0_YN3_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> CH0_YN3_ML_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          ch0_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                 // CH0_YN3_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> CH0_YN3_ML_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          ch0_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                       // CH0_YN3_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> CH0_YN3_ML_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          ch0_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;               // CH0_YN3_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> CH0_YN3_ML_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] ch0_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                        // CH0_YN3_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> CH0_YN3_ML_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          ch0_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                       // CH0_YN3_ML_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> CH0_YN3_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          ch0_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                     // CH0_YN3_ML_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> CH0_YN3_ML_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] ch0_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                      // CH0_YN3_ML_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> CH0_YN3_ML_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          ch0_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                     // CH0_YN3_ML_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> CH0_YN3_ML_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          ch0_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                           // CH0_YN3_MU_s1_translator:uav_waitrequest -> CH0_YN3_MU_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] ch0_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                            // CH0_YN3_MU_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> CH0_YN3_MU_s1_translator:uav_burstcount
	wire   [31:0] ch0_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                             // CH0_YN3_MU_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> CH0_YN3_MU_s1_translator:uav_writedata
	wire   [21:0] ch0_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_address;                               // CH0_YN3_MU_s1_translator_avalon_universal_slave_0_agent:m0_address -> CH0_YN3_MU_s1_translator:uav_address
	wire          ch0_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_write;                                 // CH0_YN3_MU_s1_translator_avalon_universal_slave_0_agent:m0_write -> CH0_YN3_MU_s1_translator:uav_write
	wire          ch0_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                  // CH0_YN3_MU_s1_translator_avalon_universal_slave_0_agent:m0_lock -> CH0_YN3_MU_s1_translator:uav_lock
	wire          ch0_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_read;                                  // CH0_YN3_MU_s1_translator_avalon_universal_slave_0_agent:m0_read -> CH0_YN3_MU_s1_translator:uav_read
	wire   [31:0] ch0_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                              // CH0_YN3_MU_s1_translator:uav_readdata -> CH0_YN3_MU_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          ch0_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                         // CH0_YN3_MU_s1_translator:uav_readdatavalid -> CH0_YN3_MU_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          ch0_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                           // CH0_YN3_MU_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> CH0_YN3_MU_s1_translator:uav_debugaccess
	wire    [3:0] ch0_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                            // CH0_YN3_MU_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> CH0_YN3_MU_s1_translator:uav_byteenable
	wire          ch0_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                    // CH0_YN3_MU_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> CH0_YN3_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          ch0_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                          // CH0_YN3_MU_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> CH0_YN3_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          ch0_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                  // CH0_YN3_MU_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> CH0_YN3_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] ch0_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                           // CH0_YN3_MU_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> CH0_YN3_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          ch0_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                          // CH0_YN3_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> CH0_YN3_MU_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          ch0_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                 // CH0_YN3_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> CH0_YN3_MU_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          ch0_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                       // CH0_YN3_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> CH0_YN3_MU_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          ch0_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;               // CH0_YN3_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> CH0_YN3_MU_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] ch0_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                        // CH0_YN3_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> CH0_YN3_MU_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          ch0_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                       // CH0_YN3_MU_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> CH0_YN3_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          ch0_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                     // CH0_YN3_MU_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> CH0_YN3_MU_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] ch0_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                      // CH0_YN3_MU_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> CH0_YN3_MU_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          ch0_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                     // CH0_YN3_MU_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> CH0_YN3_MU_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          ch0_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                            // CH0_YN3_U_s1_translator:uav_waitrequest -> CH0_YN3_U_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] ch0_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                             // CH0_YN3_U_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> CH0_YN3_U_s1_translator:uav_burstcount
	wire   [31:0] ch0_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                              // CH0_YN3_U_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> CH0_YN3_U_s1_translator:uav_writedata
	wire   [21:0] ch0_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_address;                                // CH0_YN3_U_s1_translator_avalon_universal_slave_0_agent:m0_address -> CH0_YN3_U_s1_translator:uav_address
	wire          ch0_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_write;                                  // CH0_YN3_U_s1_translator_avalon_universal_slave_0_agent:m0_write -> CH0_YN3_U_s1_translator:uav_write
	wire          ch0_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                   // CH0_YN3_U_s1_translator_avalon_universal_slave_0_agent:m0_lock -> CH0_YN3_U_s1_translator:uav_lock
	wire          ch0_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_read;                                   // CH0_YN3_U_s1_translator_avalon_universal_slave_0_agent:m0_read -> CH0_YN3_U_s1_translator:uav_read
	wire   [31:0] ch0_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                               // CH0_YN3_U_s1_translator:uav_readdata -> CH0_YN3_U_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          ch0_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                          // CH0_YN3_U_s1_translator:uav_readdatavalid -> CH0_YN3_U_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          ch0_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                            // CH0_YN3_U_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> CH0_YN3_U_s1_translator:uav_debugaccess
	wire    [3:0] ch0_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                             // CH0_YN3_U_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> CH0_YN3_U_s1_translator:uav_byteenable
	wire          ch0_yn3_u_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                     // CH0_YN3_U_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> CH0_YN3_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          ch0_yn3_u_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                           // CH0_YN3_U_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> CH0_YN3_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          ch0_yn3_u_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                   // CH0_YN3_U_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> CH0_YN3_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] ch0_yn3_u_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                            // CH0_YN3_U_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> CH0_YN3_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          ch0_yn3_u_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                           // CH0_YN3_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> CH0_YN3_U_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          ch0_yn3_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                  // CH0_YN3_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> CH0_YN3_U_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          ch0_yn3_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                        // CH0_YN3_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> CH0_YN3_U_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          ch0_yn3_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                // CH0_YN3_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> CH0_YN3_U_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] ch0_yn3_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                         // CH0_YN3_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> CH0_YN3_U_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          ch0_yn3_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                        // CH0_YN3_U_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> CH0_YN3_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          ch0_yn3_u_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                      // CH0_YN3_U_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> CH0_YN3_U_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] ch0_yn3_u_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                       // CH0_YN3_U_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> CH0_YN3_U_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          ch0_yn3_u_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                      // CH0_YN3_U_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> CH0_YN3_U_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          ch1_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                        // CH1_TIMER_RST_s1_translator:uav_waitrequest -> CH1_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] ch1_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                         // CH1_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> CH1_TIMER_RST_s1_translator:uav_burstcount
	wire   [31:0] ch1_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                          // CH1_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> CH1_TIMER_RST_s1_translator:uav_writedata
	wire   [21:0] ch1_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_address;                            // CH1_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:m0_address -> CH1_TIMER_RST_s1_translator:uav_address
	wire          ch1_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_write;                              // CH1_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:m0_write -> CH1_TIMER_RST_s1_translator:uav_write
	wire          ch1_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_lock;                               // CH1_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:m0_lock -> CH1_TIMER_RST_s1_translator:uav_lock
	wire          ch1_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_read;                               // CH1_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:m0_read -> CH1_TIMER_RST_s1_translator:uav_read
	wire   [31:0] ch1_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                           // CH1_TIMER_RST_s1_translator:uav_readdata -> CH1_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          ch1_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                      // CH1_TIMER_RST_s1_translator:uav_readdatavalid -> CH1_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          ch1_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                        // CH1_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> CH1_TIMER_RST_s1_translator:uav_debugaccess
	wire    [3:0] ch1_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                         // CH1_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> CH1_TIMER_RST_s1_translator:uav_byteenable
	wire          ch1_timer_rst_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                 // CH1_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> CH1_TIMER_RST_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          ch1_timer_rst_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                       // CH1_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> CH1_TIMER_RST_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          ch1_timer_rst_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;               // CH1_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> CH1_TIMER_RST_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] ch1_timer_rst_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                        // CH1_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> CH1_TIMER_RST_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          ch1_timer_rst_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                       // CH1_TIMER_RST_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> CH1_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          ch1_timer_rst_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;              // CH1_TIMER_RST_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> CH1_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          ch1_timer_rst_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                    // CH1_TIMER_RST_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> CH1_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          ch1_timer_rst_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;            // CH1_TIMER_RST_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> CH1_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] ch1_timer_rst_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                     // CH1_TIMER_RST_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> CH1_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          ch1_timer_rst_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                    // CH1_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> CH1_TIMER_RST_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          ch1_timer_rst_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                  // CH1_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> CH1_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] ch1_timer_rst_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                   // CH1_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> CH1_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          ch1_timer_rst_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                  // CH1_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> CH1_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          ch1_thresh_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                           // CH1_THRESH_s1_translator:uav_waitrequest -> CH1_THRESH_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] ch1_thresh_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                            // CH1_THRESH_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> CH1_THRESH_s1_translator:uav_burstcount
	wire   [31:0] ch1_thresh_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                             // CH1_THRESH_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> CH1_THRESH_s1_translator:uav_writedata
	wire   [21:0] ch1_thresh_s1_translator_avalon_universal_slave_0_agent_m0_address;                               // CH1_THRESH_s1_translator_avalon_universal_slave_0_agent:m0_address -> CH1_THRESH_s1_translator:uav_address
	wire          ch1_thresh_s1_translator_avalon_universal_slave_0_agent_m0_write;                                 // CH1_THRESH_s1_translator_avalon_universal_slave_0_agent:m0_write -> CH1_THRESH_s1_translator:uav_write
	wire          ch1_thresh_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                  // CH1_THRESH_s1_translator_avalon_universal_slave_0_agent:m0_lock -> CH1_THRESH_s1_translator:uav_lock
	wire          ch1_thresh_s1_translator_avalon_universal_slave_0_agent_m0_read;                                  // CH1_THRESH_s1_translator_avalon_universal_slave_0_agent:m0_read -> CH1_THRESH_s1_translator:uav_read
	wire   [31:0] ch1_thresh_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                              // CH1_THRESH_s1_translator:uav_readdata -> CH1_THRESH_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          ch1_thresh_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                         // CH1_THRESH_s1_translator:uav_readdatavalid -> CH1_THRESH_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          ch1_thresh_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                           // CH1_THRESH_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> CH1_THRESH_s1_translator:uav_debugaccess
	wire    [3:0] ch1_thresh_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                            // CH1_THRESH_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> CH1_THRESH_s1_translator:uav_byteenable
	wire          ch1_thresh_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                    // CH1_THRESH_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> CH1_THRESH_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          ch1_thresh_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                          // CH1_THRESH_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> CH1_THRESH_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          ch1_thresh_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                  // CH1_THRESH_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> CH1_THRESH_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] ch1_thresh_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                           // CH1_THRESH_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> CH1_THRESH_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          ch1_thresh_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                          // CH1_THRESH_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> CH1_THRESH_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          ch1_thresh_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                 // CH1_THRESH_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> CH1_THRESH_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          ch1_thresh_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                       // CH1_THRESH_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> CH1_THRESH_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          ch1_thresh_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;               // CH1_THRESH_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> CH1_THRESH_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] ch1_thresh_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                        // CH1_THRESH_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> CH1_THRESH_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          ch1_thresh_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                       // CH1_THRESH_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> CH1_THRESH_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          ch1_thresh_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                     // CH1_THRESH_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> CH1_THRESH_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] ch1_thresh_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                      // CH1_THRESH_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> CH1_THRESH_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          ch1_thresh_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                     // CH1_THRESH_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> CH1_THRESH_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          ch1_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                          // CH1_RD_PEAK_s1_translator:uav_waitrequest -> CH1_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] ch1_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                           // CH1_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> CH1_RD_PEAK_s1_translator:uav_burstcount
	wire   [31:0] ch1_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                            // CH1_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> CH1_RD_PEAK_s1_translator:uav_writedata
	wire   [21:0] ch1_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_address;                              // CH1_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:m0_address -> CH1_RD_PEAK_s1_translator:uav_address
	wire          ch1_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_write;                                // CH1_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:m0_write -> CH1_RD_PEAK_s1_translator:uav_write
	wire          ch1_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                 // CH1_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:m0_lock -> CH1_RD_PEAK_s1_translator:uav_lock
	wire          ch1_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_read;                                 // CH1_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:m0_read -> CH1_RD_PEAK_s1_translator:uav_read
	wire   [31:0] ch1_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                             // CH1_RD_PEAK_s1_translator:uav_readdata -> CH1_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          ch1_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                        // CH1_RD_PEAK_s1_translator:uav_readdatavalid -> CH1_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          ch1_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                          // CH1_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> CH1_RD_PEAK_s1_translator:uav_debugaccess
	wire    [3:0] ch1_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                           // CH1_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> CH1_RD_PEAK_s1_translator:uav_byteenable
	wire          ch1_rd_peak_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                   // CH1_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> CH1_RD_PEAK_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          ch1_rd_peak_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                         // CH1_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> CH1_RD_PEAK_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          ch1_rd_peak_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                 // CH1_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> CH1_RD_PEAK_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] ch1_rd_peak_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                          // CH1_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> CH1_RD_PEAK_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          ch1_rd_peak_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                         // CH1_RD_PEAK_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> CH1_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          ch1_rd_peak_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                // CH1_RD_PEAK_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> CH1_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          ch1_rd_peak_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                      // CH1_RD_PEAK_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> CH1_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          ch1_rd_peak_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;              // CH1_RD_PEAK_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> CH1_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] ch1_rd_peak_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                       // CH1_RD_PEAK_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> CH1_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          ch1_rd_peak_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                      // CH1_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> CH1_RD_PEAK_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          ch1_rd_peak_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                    // CH1_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> CH1_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] ch1_rd_peak_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                     // CH1_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> CH1_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          ch1_rd_peak_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                    // CH1_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> CH1_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          ch1_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                       // CH1_PEAK_FOUND_s1_translator:uav_waitrequest -> CH1_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] ch1_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                        // CH1_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> CH1_PEAK_FOUND_s1_translator:uav_burstcount
	wire   [31:0] ch1_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                         // CH1_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> CH1_PEAK_FOUND_s1_translator:uav_writedata
	wire   [21:0] ch1_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_address;                           // CH1_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:m0_address -> CH1_PEAK_FOUND_s1_translator:uav_address
	wire          ch1_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_write;                             // CH1_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:m0_write -> CH1_PEAK_FOUND_s1_translator:uav_write
	wire          ch1_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_lock;                              // CH1_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:m0_lock -> CH1_PEAK_FOUND_s1_translator:uav_lock
	wire          ch1_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_read;                              // CH1_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:m0_read -> CH1_PEAK_FOUND_s1_translator:uav_read
	wire   [31:0] ch1_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                          // CH1_PEAK_FOUND_s1_translator:uav_readdata -> CH1_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          ch1_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                     // CH1_PEAK_FOUND_s1_translator:uav_readdatavalid -> CH1_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          ch1_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                       // CH1_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> CH1_PEAK_FOUND_s1_translator:uav_debugaccess
	wire    [3:0] ch1_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                        // CH1_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> CH1_PEAK_FOUND_s1_translator:uav_byteenable
	wire          ch1_peak_found_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                // CH1_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> CH1_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          ch1_peak_found_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                      // CH1_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> CH1_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          ch1_peak_found_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;              // CH1_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> CH1_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] ch1_peak_found_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                       // CH1_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> CH1_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          ch1_peak_found_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                      // CH1_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> CH1_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          ch1_peak_found_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;             // CH1_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> CH1_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          ch1_peak_found_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                   // CH1_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> CH1_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          ch1_peak_found_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;           // CH1_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> CH1_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] ch1_peak_found_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                    // CH1_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> CH1_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          ch1_peak_found_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                   // CH1_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> CH1_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          ch1_peak_found_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                 // CH1_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> CH1_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] ch1_peak_found_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                  // CH1_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> CH1_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          ch1_peak_found_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                 // CH1_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> CH1_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          ch1_time_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                             // CH1_TIME_s1_translator:uav_waitrequest -> CH1_TIME_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] ch1_time_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                              // CH1_TIME_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> CH1_TIME_s1_translator:uav_burstcount
	wire   [31:0] ch1_time_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                               // CH1_TIME_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> CH1_TIME_s1_translator:uav_writedata
	wire   [21:0] ch1_time_s1_translator_avalon_universal_slave_0_agent_m0_address;                                 // CH1_TIME_s1_translator_avalon_universal_slave_0_agent:m0_address -> CH1_TIME_s1_translator:uav_address
	wire          ch1_time_s1_translator_avalon_universal_slave_0_agent_m0_write;                                   // CH1_TIME_s1_translator_avalon_universal_slave_0_agent:m0_write -> CH1_TIME_s1_translator:uav_write
	wire          ch1_time_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                    // CH1_TIME_s1_translator_avalon_universal_slave_0_agent:m0_lock -> CH1_TIME_s1_translator:uav_lock
	wire          ch1_time_s1_translator_avalon_universal_slave_0_agent_m0_read;                                    // CH1_TIME_s1_translator_avalon_universal_slave_0_agent:m0_read -> CH1_TIME_s1_translator:uav_read
	wire   [31:0] ch1_time_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                // CH1_TIME_s1_translator:uav_readdata -> CH1_TIME_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          ch1_time_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                           // CH1_TIME_s1_translator:uav_readdatavalid -> CH1_TIME_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          ch1_time_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                             // CH1_TIME_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> CH1_TIME_s1_translator:uav_debugaccess
	wire    [3:0] ch1_time_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                              // CH1_TIME_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> CH1_TIME_s1_translator:uav_byteenable
	wire          ch1_time_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                      // CH1_TIME_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> CH1_TIME_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          ch1_time_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                            // CH1_TIME_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> CH1_TIME_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          ch1_time_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                    // CH1_TIME_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> CH1_TIME_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] ch1_time_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                             // CH1_TIME_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> CH1_TIME_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          ch1_time_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                            // CH1_TIME_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> CH1_TIME_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          ch1_time_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                   // CH1_TIME_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> CH1_TIME_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          ch1_time_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                         // CH1_TIME_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> CH1_TIME_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          ch1_time_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                 // CH1_TIME_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> CH1_TIME_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] ch1_time_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                          // CH1_TIME_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> CH1_TIME_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          ch1_time_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                         // CH1_TIME_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> CH1_TIME_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          ch1_time_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                       // CH1_TIME_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> CH1_TIME_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] ch1_time_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                        // CH1_TIME_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> CH1_TIME_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          ch1_time_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                       // CH1_TIME_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> CH1_TIME_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          ch1_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                            // CH1_YN1_U_s1_translator:uav_waitrequest -> CH1_YN1_U_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] ch1_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                             // CH1_YN1_U_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> CH1_YN1_U_s1_translator:uav_burstcount
	wire   [31:0] ch1_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                              // CH1_YN1_U_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> CH1_YN1_U_s1_translator:uav_writedata
	wire   [21:0] ch1_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_address;                                // CH1_YN1_U_s1_translator_avalon_universal_slave_0_agent:m0_address -> CH1_YN1_U_s1_translator:uav_address
	wire          ch1_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_write;                                  // CH1_YN1_U_s1_translator_avalon_universal_slave_0_agent:m0_write -> CH1_YN1_U_s1_translator:uav_write
	wire          ch1_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                   // CH1_YN1_U_s1_translator_avalon_universal_slave_0_agent:m0_lock -> CH1_YN1_U_s1_translator:uav_lock
	wire          ch1_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_read;                                   // CH1_YN1_U_s1_translator_avalon_universal_slave_0_agent:m0_read -> CH1_YN1_U_s1_translator:uav_read
	wire   [31:0] ch1_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                               // CH1_YN1_U_s1_translator:uav_readdata -> CH1_YN1_U_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          ch1_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                          // CH1_YN1_U_s1_translator:uav_readdatavalid -> CH1_YN1_U_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          ch1_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                            // CH1_YN1_U_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> CH1_YN1_U_s1_translator:uav_debugaccess
	wire    [3:0] ch1_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                             // CH1_YN1_U_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> CH1_YN1_U_s1_translator:uav_byteenable
	wire          ch1_yn1_u_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                     // CH1_YN1_U_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> CH1_YN1_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          ch1_yn1_u_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                           // CH1_YN1_U_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> CH1_YN1_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          ch1_yn1_u_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                   // CH1_YN1_U_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> CH1_YN1_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] ch1_yn1_u_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                            // CH1_YN1_U_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> CH1_YN1_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          ch1_yn1_u_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                           // CH1_YN1_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> CH1_YN1_U_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          ch1_yn1_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                  // CH1_YN1_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> CH1_YN1_U_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          ch1_yn1_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                        // CH1_YN1_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> CH1_YN1_U_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          ch1_yn1_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                // CH1_YN1_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> CH1_YN1_U_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] ch1_yn1_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                         // CH1_YN1_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> CH1_YN1_U_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          ch1_yn1_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                        // CH1_YN1_U_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> CH1_YN1_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          ch1_yn1_u_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                      // CH1_YN1_U_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> CH1_YN1_U_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] ch1_yn1_u_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                       // CH1_YN1_U_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> CH1_YN1_U_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          ch1_yn1_u_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                      // CH1_YN1_U_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> CH1_YN1_U_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          ch1_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                           // CH1_YN1_MU_s1_translator:uav_waitrequest -> CH1_YN1_MU_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] ch1_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                            // CH1_YN1_MU_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> CH1_YN1_MU_s1_translator:uav_burstcount
	wire   [31:0] ch1_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                             // CH1_YN1_MU_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> CH1_YN1_MU_s1_translator:uav_writedata
	wire   [21:0] ch1_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_address;                               // CH1_YN1_MU_s1_translator_avalon_universal_slave_0_agent:m0_address -> CH1_YN1_MU_s1_translator:uav_address
	wire          ch1_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_write;                                 // CH1_YN1_MU_s1_translator_avalon_universal_slave_0_agent:m0_write -> CH1_YN1_MU_s1_translator:uav_write
	wire          ch1_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                  // CH1_YN1_MU_s1_translator_avalon_universal_slave_0_agent:m0_lock -> CH1_YN1_MU_s1_translator:uav_lock
	wire          ch1_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_read;                                  // CH1_YN1_MU_s1_translator_avalon_universal_slave_0_agent:m0_read -> CH1_YN1_MU_s1_translator:uav_read
	wire   [31:0] ch1_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                              // CH1_YN1_MU_s1_translator:uav_readdata -> CH1_YN1_MU_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          ch1_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                         // CH1_YN1_MU_s1_translator:uav_readdatavalid -> CH1_YN1_MU_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          ch1_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                           // CH1_YN1_MU_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> CH1_YN1_MU_s1_translator:uav_debugaccess
	wire    [3:0] ch1_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                            // CH1_YN1_MU_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> CH1_YN1_MU_s1_translator:uav_byteenable
	wire          ch1_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                    // CH1_YN1_MU_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> CH1_YN1_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          ch1_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                          // CH1_YN1_MU_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> CH1_YN1_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          ch1_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                  // CH1_YN1_MU_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> CH1_YN1_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] ch1_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                           // CH1_YN1_MU_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> CH1_YN1_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          ch1_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                          // CH1_YN1_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> CH1_YN1_MU_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          ch1_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                 // CH1_YN1_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> CH1_YN1_MU_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          ch1_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                       // CH1_YN1_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> CH1_YN1_MU_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          ch1_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;               // CH1_YN1_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> CH1_YN1_MU_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] ch1_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                        // CH1_YN1_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> CH1_YN1_MU_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          ch1_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                       // CH1_YN1_MU_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> CH1_YN1_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          ch1_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                     // CH1_YN1_MU_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> CH1_YN1_MU_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] ch1_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                      // CH1_YN1_MU_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> CH1_YN1_MU_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          ch1_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                     // CH1_YN1_MU_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> CH1_YN1_MU_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          ch1_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                           // CH1_YN1_ML_s1_translator:uav_waitrequest -> CH1_YN1_ML_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] ch1_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                            // CH1_YN1_ML_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> CH1_YN1_ML_s1_translator:uav_burstcount
	wire   [31:0] ch1_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                             // CH1_YN1_ML_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> CH1_YN1_ML_s1_translator:uav_writedata
	wire   [21:0] ch1_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_address;                               // CH1_YN1_ML_s1_translator_avalon_universal_slave_0_agent:m0_address -> CH1_YN1_ML_s1_translator:uav_address
	wire          ch1_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_write;                                 // CH1_YN1_ML_s1_translator_avalon_universal_slave_0_agent:m0_write -> CH1_YN1_ML_s1_translator:uav_write
	wire          ch1_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                  // CH1_YN1_ML_s1_translator_avalon_universal_slave_0_agent:m0_lock -> CH1_YN1_ML_s1_translator:uav_lock
	wire          ch1_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_read;                                  // CH1_YN1_ML_s1_translator_avalon_universal_slave_0_agent:m0_read -> CH1_YN1_ML_s1_translator:uav_read
	wire   [31:0] ch1_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                              // CH1_YN1_ML_s1_translator:uav_readdata -> CH1_YN1_ML_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          ch1_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                         // CH1_YN1_ML_s1_translator:uav_readdatavalid -> CH1_YN1_ML_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          ch1_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                           // CH1_YN1_ML_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> CH1_YN1_ML_s1_translator:uav_debugaccess
	wire    [3:0] ch1_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                            // CH1_YN1_ML_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> CH1_YN1_ML_s1_translator:uav_byteenable
	wire          ch1_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                    // CH1_YN1_ML_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> CH1_YN1_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          ch1_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                          // CH1_YN1_ML_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> CH1_YN1_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          ch1_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                  // CH1_YN1_ML_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> CH1_YN1_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] ch1_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                           // CH1_YN1_ML_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> CH1_YN1_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          ch1_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                          // CH1_YN1_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> CH1_YN1_ML_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          ch1_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                 // CH1_YN1_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> CH1_YN1_ML_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          ch1_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                       // CH1_YN1_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> CH1_YN1_ML_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          ch1_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;               // CH1_YN1_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> CH1_YN1_ML_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] ch1_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                        // CH1_YN1_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> CH1_YN1_ML_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          ch1_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                       // CH1_YN1_ML_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> CH1_YN1_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          ch1_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                     // CH1_YN1_ML_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> CH1_YN1_ML_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] ch1_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                      // CH1_YN1_ML_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> CH1_YN1_ML_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          ch1_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                     // CH1_YN1_ML_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> CH1_YN1_ML_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          ch1_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                            // CH1_YN1_L_s1_translator:uav_waitrequest -> CH1_YN1_L_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] ch1_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                             // CH1_YN1_L_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> CH1_YN1_L_s1_translator:uav_burstcount
	wire   [31:0] ch1_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                              // CH1_YN1_L_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> CH1_YN1_L_s1_translator:uav_writedata
	wire   [21:0] ch1_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_address;                                // CH1_YN1_L_s1_translator_avalon_universal_slave_0_agent:m0_address -> CH1_YN1_L_s1_translator:uav_address
	wire          ch1_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_write;                                  // CH1_YN1_L_s1_translator_avalon_universal_slave_0_agent:m0_write -> CH1_YN1_L_s1_translator:uav_write
	wire          ch1_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                   // CH1_YN1_L_s1_translator_avalon_universal_slave_0_agent:m0_lock -> CH1_YN1_L_s1_translator:uav_lock
	wire          ch1_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_read;                                   // CH1_YN1_L_s1_translator_avalon_universal_slave_0_agent:m0_read -> CH1_YN1_L_s1_translator:uav_read
	wire   [31:0] ch1_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                               // CH1_YN1_L_s1_translator:uav_readdata -> CH1_YN1_L_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          ch1_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                          // CH1_YN1_L_s1_translator:uav_readdatavalid -> CH1_YN1_L_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          ch1_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                            // CH1_YN1_L_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> CH1_YN1_L_s1_translator:uav_debugaccess
	wire    [3:0] ch1_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                             // CH1_YN1_L_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> CH1_YN1_L_s1_translator:uav_byteenable
	wire          ch1_yn1_l_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                     // CH1_YN1_L_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> CH1_YN1_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          ch1_yn1_l_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                           // CH1_YN1_L_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> CH1_YN1_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          ch1_yn1_l_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                   // CH1_YN1_L_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> CH1_YN1_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] ch1_yn1_l_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                            // CH1_YN1_L_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> CH1_YN1_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          ch1_yn1_l_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                           // CH1_YN1_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> CH1_YN1_L_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          ch1_yn1_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                  // CH1_YN1_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> CH1_YN1_L_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          ch1_yn1_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                        // CH1_YN1_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> CH1_YN1_L_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          ch1_yn1_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                // CH1_YN1_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> CH1_YN1_L_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] ch1_yn1_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                         // CH1_YN1_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> CH1_YN1_L_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          ch1_yn1_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                        // CH1_YN1_L_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> CH1_YN1_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          ch1_yn1_l_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                      // CH1_YN1_L_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> CH1_YN1_L_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] ch1_yn1_l_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                       // CH1_YN1_L_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> CH1_YN1_L_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          ch1_yn1_l_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                      // CH1_YN1_L_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> CH1_YN1_L_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          ch1_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                            // CH1_YN2_U_s1_translator:uav_waitrequest -> CH1_YN2_U_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] ch1_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                             // CH1_YN2_U_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> CH1_YN2_U_s1_translator:uav_burstcount
	wire   [31:0] ch1_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                              // CH1_YN2_U_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> CH1_YN2_U_s1_translator:uav_writedata
	wire   [21:0] ch1_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_address;                                // CH1_YN2_U_s1_translator_avalon_universal_slave_0_agent:m0_address -> CH1_YN2_U_s1_translator:uav_address
	wire          ch1_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_write;                                  // CH1_YN2_U_s1_translator_avalon_universal_slave_0_agent:m0_write -> CH1_YN2_U_s1_translator:uav_write
	wire          ch1_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                   // CH1_YN2_U_s1_translator_avalon_universal_slave_0_agent:m0_lock -> CH1_YN2_U_s1_translator:uav_lock
	wire          ch1_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_read;                                   // CH1_YN2_U_s1_translator_avalon_universal_slave_0_agent:m0_read -> CH1_YN2_U_s1_translator:uav_read
	wire   [31:0] ch1_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                               // CH1_YN2_U_s1_translator:uav_readdata -> CH1_YN2_U_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          ch1_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                          // CH1_YN2_U_s1_translator:uav_readdatavalid -> CH1_YN2_U_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          ch1_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                            // CH1_YN2_U_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> CH1_YN2_U_s1_translator:uav_debugaccess
	wire    [3:0] ch1_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                             // CH1_YN2_U_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> CH1_YN2_U_s1_translator:uav_byteenable
	wire          ch1_yn2_u_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                     // CH1_YN2_U_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> CH1_YN2_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          ch1_yn2_u_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                           // CH1_YN2_U_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> CH1_YN2_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          ch1_yn2_u_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                   // CH1_YN2_U_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> CH1_YN2_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] ch1_yn2_u_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                            // CH1_YN2_U_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> CH1_YN2_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          ch1_yn2_u_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                           // CH1_YN2_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> CH1_YN2_U_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          ch1_yn2_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                  // CH1_YN2_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> CH1_YN2_U_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          ch1_yn2_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                        // CH1_YN2_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> CH1_YN2_U_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          ch1_yn2_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                // CH1_YN2_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> CH1_YN2_U_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] ch1_yn2_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                         // CH1_YN2_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> CH1_YN2_U_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          ch1_yn2_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                        // CH1_YN2_U_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> CH1_YN2_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          ch1_yn2_u_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                      // CH1_YN2_U_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> CH1_YN2_U_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] ch1_yn2_u_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                       // CH1_YN2_U_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> CH1_YN2_U_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          ch1_yn2_u_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                      // CH1_YN2_U_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> CH1_YN2_U_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          ch1_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                           // CH1_YN2_MU_s1_translator:uav_waitrequest -> CH1_YN2_MU_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] ch1_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                            // CH1_YN2_MU_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> CH1_YN2_MU_s1_translator:uav_burstcount
	wire   [31:0] ch1_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                             // CH1_YN2_MU_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> CH1_YN2_MU_s1_translator:uav_writedata
	wire   [21:0] ch1_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_address;                               // CH1_YN2_MU_s1_translator_avalon_universal_slave_0_agent:m0_address -> CH1_YN2_MU_s1_translator:uav_address
	wire          ch1_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_write;                                 // CH1_YN2_MU_s1_translator_avalon_universal_slave_0_agent:m0_write -> CH1_YN2_MU_s1_translator:uav_write
	wire          ch1_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                  // CH1_YN2_MU_s1_translator_avalon_universal_slave_0_agent:m0_lock -> CH1_YN2_MU_s1_translator:uav_lock
	wire          ch1_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_read;                                  // CH1_YN2_MU_s1_translator_avalon_universal_slave_0_agent:m0_read -> CH1_YN2_MU_s1_translator:uav_read
	wire   [31:0] ch1_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                              // CH1_YN2_MU_s1_translator:uav_readdata -> CH1_YN2_MU_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          ch1_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                         // CH1_YN2_MU_s1_translator:uav_readdatavalid -> CH1_YN2_MU_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          ch1_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                           // CH1_YN2_MU_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> CH1_YN2_MU_s1_translator:uav_debugaccess
	wire    [3:0] ch1_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                            // CH1_YN2_MU_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> CH1_YN2_MU_s1_translator:uav_byteenable
	wire          ch1_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                    // CH1_YN2_MU_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> CH1_YN2_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          ch1_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                          // CH1_YN2_MU_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> CH1_YN2_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          ch1_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                  // CH1_YN2_MU_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> CH1_YN2_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] ch1_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                           // CH1_YN2_MU_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> CH1_YN2_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          ch1_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                          // CH1_YN2_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> CH1_YN2_MU_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          ch1_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                 // CH1_YN2_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> CH1_YN2_MU_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          ch1_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                       // CH1_YN2_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> CH1_YN2_MU_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          ch1_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;               // CH1_YN2_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> CH1_YN2_MU_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] ch1_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                        // CH1_YN2_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> CH1_YN2_MU_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          ch1_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                       // CH1_YN2_MU_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> CH1_YN2_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          ch1_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                     // CH1_YN2_MU_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> CH1_YN2_MU_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] ch1_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                      // CH1_YN2_MU_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> CH1_YN2_MU_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          ch1_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                     // CH1_YN2_MU_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> CH1_YN2_MU_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          ch1_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                           // CH1_YN2_ML_s1_translator:uav_waitrequest -> CH1_YN2_ML_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] ch1_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                            // CH1_YN2_ML_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> CH1_YN2_ML_s1_translator:uav_burstcount
	wire   [31:0] ch1_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                             // CH1_YN2_ML_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> CH1_YN2_ML_s1_translator:uav_writedata
	wire   [21:0] ch1_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_address;                               // CH1_YN2_ML_s1_translator_avalon_universal_slave_0_agent:m0_address -> CH1_YN2_ML_s1_translator:uav_address
	wire          ch1_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_write;                                 // CH1_YN2_ML_s1_translator_avalon_universal_slave_0_agent:m0_write -> CH1_YN2_ML_s1_translator:uav_write
	wire          ch1_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                  // CH1_YN2_ML_s1_translator_avalon_universal_slave_0_agent:m0_lock -> CH1_YN2_ML_s1_translator:uav_lock
	wire          ch1_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_read;                                  // CH1_YN2_ML_s1_translator_avalon_universal_slave_0_agent:m0_read -> CH1_YN2_ML_s1_translator:uav_read
	wire   [31:0] ch1_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                              // CH1_YN2_ML_s1_translator:uav_readdata -> CH1_YN2_ML_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          ch1_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                         // CH1_YN2_ML_s1_translator:uav_readdatavalid -> CH1_YN2_ML_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          ch1_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                           // CH1_YN2_ML_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> CH1_YN2_ML_s1_translator:uav_debugaccess
	wire    [3:0] ch1_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                            // CH1_YN2_ML_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> CH1_YN2_ML_s1_translator:uav_byteenable
	wire          ch1_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                    // CH1_YN2_ML_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> CH1_YN2_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          ch1_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                          // CH1_YN2_ML_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> CH1_YN2_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          ch1_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                  // CH1_YN2_ML_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> CH1_YN2_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] ch1_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                           // CH1_YN2_ML_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> CH1_YN2_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          ch1_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                          // CH1_YN2_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> CH1_YN2_ML_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          ch1_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                 // CH1_YN2_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> CH1_YN2_ML_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          ch1_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                       // CH1_YN2_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> CH1_YN2_ML_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          ch1_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;               // CH1_YN2_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> CH1_YN2_ML_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] ch1_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                        // CH1_YN2_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> CH1_YN2_ML_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          ch1_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                       // CH1_YN2_ML_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> CH1_YN2_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          ch1_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                     // CH1_YN2_ML_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> CH1_YN2_ML_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] ch1_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                      // CH1_YN2_ML_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> CH1_YN2_ML_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          ch1_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                     // CH1_YN2_ML_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> CH1_YN2_ML_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          ch1_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                            // CH1_YN2_L_s1_translator:uav_waitrequest -> CH1_YN2_L_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] ch1_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                             // CH1_YN2_L_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> CH1_YN2_L_s1_translator:uav_burstcount
	wire   [31:0] ch1_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                              // CH1_YN2_L_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> CH1_YN2_L_s1_translator:uav_writedata
	wire   [21:0] ch1_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_address;                                // CH1_YN2_L_s1_translator_avalon_universal_slave_0_agent:m0_address -> CH1_YN2_L_s1_translator:uav_address
	wire          ch1_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_write;                                  // CH1_YN2_L_s1_translator_avalon_universal_slave_0_agent:m0_write -> CH1_YN2_L_s1_translator:uav_write
	wire          ch1_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                   // CH1_YN2_L_s1_translator_avalon_universal_slave_0_agent:m0_lock -> CH1_YN2_L_s1_translator:uav_lock
	wire          ch1_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_read;                                   // CH1_YN2_L_s1_translator_avalon_universal_slave_0_agent:m0_read -> CH1_YN2_L_s1_translator:uav_read
	wire   [31:0] ch1_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                               // CH1_YN2_L_s1_translator:uav_readdata -> CH1_YN2_L_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          ch1_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                          // CH1_YN2_L_s1_translator:uav_readdatavalid -> CH1_YN2_L_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          ch1_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                            // CH1_YN2_L_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> CH1_YN2_L_s1_translator:uav_debugaccess
	wire    [3:0] ch1_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                             // CH1_YN2_L_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> CH1_YN2_L_s1_translator:uav_byteenable
	wire          ch1_yn2_l_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                     // CH1_YN2_L_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> CH1_YN2_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          ch1_yn2_l_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                           // CH1_YN2_L_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> CH1_YN2_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          ch1_yn2_l_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                   // CH1_YN2_L_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> CH1_YN2_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] ch1_yn2_l_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                            // CH1_YN2_L_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> CH1_YN2_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          ch1_yn2_l_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                           // CH1_YN2_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> CH1_YN2_L_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          ch1_yn2_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                  // CH1_YN2_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> CH1_YN2_L_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          ch1_yn2_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                        // CH1_YN2_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> CH1_YN2_L_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          ch1_yn2_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                // CH1_YN2_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> CH1_YN2_L_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] ch1_yn2_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                         // CH1_YN2_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> CH1_YN2_L_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          ch1_yn2_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                        // CH1_YN2_L_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> CH1_YN2_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          ch1_yn2_l_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                      // CH1_YN2_L_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> CH1_YN2_L_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] ch1_yn2_l_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                       // CH1_YN2_L_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> CH1_YN2_L_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          ch1_yn2_l_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                      // CH1_YN2_L_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> CH1_YN2_L_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          ch1_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                            // CH1_YN3_U_s1_translator:uav_waitrequest -> CH1_YN3_U_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] ch1_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                             // CH1_YN3_U_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> CH1_YN3_U_s1_translator:uav_burstcount
	wire   [31:0] ch1_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                              // CH1_YN3_U_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> CH1_YN3_U_s1_translator:uav_writedata
	wire   [21:0] ch1_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_address;                                // CH1_YN3_U_s1_translator_avalon_universal_slave_0_agent:m0_address -> CH1_YN3_U_s1_translator:uav_address
	wire          ch1_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_write;                                  // CH1_YN3_U_s1_translator_avalon_universal_slave_0_agent:m0_write -> CH1_YN3_U_s1_translator:uav_write
	wire          ch1_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                   // CH1_YN3_U_s1_translator_avalon_universal_slave_0_agent:m0_lock -> CH1_YN3_U_s1_translator:uav_lock
	wire          ch1_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_read;                                   // CH1_YN3_U_s1_translator_avalon_universal_slave_0_agent:m0_read -> CH1_YN3_U_s1_translator:uav_read
	wire   [31:0] ch1_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                               // CH1_YN3_U_s1_translator:uav_readdata -> CH1_YN3_U_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          ch1_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                          // CH1_YN3_U_s1_translator:uav_readdatavalid -> CH1_YN3_U_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          ch1_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                            // CH1_YN3_U_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> CH1_YN3_U_s1_translator:uav_debugaccess
	wire    [3:0] ch1_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                             // CH1_YN3_U_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> CH1_YN3_U_s1_translator:uav_byteenable
	wire          ch1_yn3_u_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                     // CH1_YN3_U_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> CH1_YN3_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          ch1_yn3_u_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                           // CH1_YN3_U_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> CH1_YN3_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          ch1_yn3_u_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                   // CH1_YN3_U_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> CH1_YN3_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] ch1_yn3_u_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                            // CH1_YN3_U_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> CH1_YN3_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          ch1_yn3_u_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                           // CH1_YN3_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> CH1_YN3_U_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          ch1_yn3_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                  // CH1_YN3_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> CH1_YN3_U_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          ch1_yn3_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                        // CH1_YN3_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> CH1_YN3_U_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          ch1_yn3_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                // CH1_YN3_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> CH1_YN3_U_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] ch1_yn3_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                         // CH1_YN3_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> CH1_YN3_U_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          ch1_yn3_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                        // CH1_YN3_U_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> CH1_YN3_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          ch1_yn3_u_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                      // CH1_YN3_U_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> CH1_YN3_U_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] ch1_yn3_u_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                       // CH1_YN3_U_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> CH1_YN3_U_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          ch1_yn3_u_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                      // CH1_YN3_U_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> CH1_YN3_U_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          ch1_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                           // CH1_YN3_MU_s1_translator:uav_waitrequest -> CH1_YN3_MU_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] ch1_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                            // CH1_YN3_MU_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> CH1_YN3_MU_s1_translator:uav_burstcount
	wire   [31:0] ch1_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                             // CH1_YN3_MU_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> CH1_YN3_MU_s1_translator:uav_writedata
	wire   [21:0] ch1_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_address;                               // CH1_YN3_MU_s1_translator_avalon_universal_slave_0_agent:m0_address -> CH1_YN3_MU_s1_translator:uav_address
	wire          ch1_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_write;                                 // CH1_YN3_MU_s1_translator_avalon_universal_slave_0_agent:m0_write -> CH1_YN3_MU_s1_translator:uav_write
	wire          ch1_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                  // CH1_YN3_MU_s1_translator_avalon_universal_slave_0_agent:m0_lock -> CH1_YN3_MU_s1_translator:uav_lock
	wire          ch1_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_read;                                  // CH1_YN3_MU_s1_translator_avalon_universal_slave_0_agent:m0_read -> CH1_YN3_MU_s1_translator:uav_read
	wire   [31:0] ch1_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                              // CH1_YN3_MU_s1_translator:uav_readdata -> CH1_YN3_MU_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          ch1_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                         // CH1_YN3_MU_s1_translator:uav_readdatavalid -> CH1_YN3_MU_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          ch1_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                           // CH1_YN3_MU_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> CH1_YN3_MU_s1_translator:uav_debugaccess
	wire    [3:0] ch1_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                            // CH1_YN3_MU_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> CH1_YN3_MU_s1_translator:uav_byteenable
	wire          ch1_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                    // CH1_YN3_MU_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> CH1_YN3_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          ch1_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                          // CH1_YN3_MU_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> CH1_YN3_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          ch1_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                  // CH1_YN3_MU_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> CH1_YN3_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] ch1_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                           // CH1_YN3_MU_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> CH1_YN3_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          ch1_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                          // CH1_YN3_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> CH1_YN3_MU_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          ch1_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                 // CH1_YN3_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> CH1_YN3_MU_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          ch1_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                       // CH1_YN3_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> CH1_YN3_MU_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          ch1_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;               // CH1_YN3_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> CH1_YN3_MU_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] ch1_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                        // CH1_YN3_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> CH1_YN3_MU_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          ch1_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                       // CH1_YN3_MU_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> CH1_YN3_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          ch1_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                     // CH1_YN3_MU_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> CH1_YN3_MU_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] ch1_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                      // CH1_YN3_MU_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> CH1_YN3_MU_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          ch1_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                     // CH1_YN3_MU_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> CH1_YN3_MU_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          ch1_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                           // CH1_YN3_ML_s1_translator:uav_waitrequest -> CH1_YN3_ML_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] ch1_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                            // CH1_YN3_ML_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> CH1_YN3_ML_s1_translator:uav_burstcount
	wire   [31:0] ch1_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                             // CH1_YN3_ML_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> CH1_YN3_ML_s1_translator:uav_writedata
	wire   [21:0] ch1_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_address;                               // CH1_YN3_ML_s1_translator_avalon_universal_slave_0_agent:m0_address -> CH1_YN3_ML_s1_translator:uav_address
	wire          ch1_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_write;                                 // CH1_YN3_ML_s1_translator_avalon_universal_slave_0_agent:m0_write -> CH1_YN3_ML_s1_translator:uav_write
	wire          ch1_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                  // CH1_YN3_ML_s1_translator_avalon_universal_slave_0_agent:m0_lock -> CH1_YN3_ML_s1_translator:uav_lock
	wire          ch1_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_read;                                  // CH1_YN3_ML_s1_translator_avalon_universal_slave_0_agent:m0_read -> CH1_YN3_ML_s1_translator:uav_read
	wire   [31:0] ch1_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                              // CH1_YN3_ML_s1_translator:uav_readdata -> CH1_YN3_ML_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          ch1_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                         // CH1_YN3_ML_s1_translator:uav_readdatavalid -> CH1_YN3_ML_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          ch1_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                           // CH1_YN3_ML_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> CH1_YN3_ML_s1_translator:uav_debugaccess
	wire    [3:0] ch1_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                            // CH1_YN3_ML_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> CH1_YN3_ML_s1_translator:uav_byteenable
	wire          ch1_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                    // CH1_YN3_ML_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> CH1_YN3_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          ch1_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                          // CH1_YN3_ML_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> CH1_YN3_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          ch1_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                  // CH1_YN3_ML_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> CH1_YN3_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] ch1_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                           // CH1_YN3_ML_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> CH1_YN3_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          ch1_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                          // CH1_YN3_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> CH1_YN3_ML_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          ch1_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                 // CH1_YN3_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> CH1_YN3_ML_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          ch1_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                       // CH1_YN3_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> CH1_YN3_ML_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          ch1_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;               // CH1_YN3_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> CH1_YN3_ML_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] ch1_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                        // CH1_YN3_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> CH1_YN3_ML_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          ch1_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                       // CH1_YN3_ML_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> CH1_YN3_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          ch1_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                     // CH1_YN3_ML_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> CH1_YN3_ML_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] ch1_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                      // CH1_YN3_ML_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> CH1_YN3_ML_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          ch1_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                     // CH1_YN3_ML_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> CH1_YN3_ML_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          ch1_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                            // CH1_YN3_L_s1_translator:uav_waitrequest -> CH1_YN3_L_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] ch1_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                             // CH1_YN3_L_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> CH1_YN3_L_s1_translator:uav_burstcount
	wire   [31:0] ch1_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                              // CH1_YN3_L_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> CH1_YN3_L_s1_translator:uav_writedata
	wire   [21:0] ch1_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_address;                                // CH1_YN3_L_s1_translator_avalon_universal_slave_0_agent:m0_address -> CH1_YN3_L_s1_translator:uav_address
	wire          ch1_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_write;                                  // CH1_YN3_L_s1_translator_avalon_universal_slave_0_agent:m0_write -> CH1_YN3_L_s1_translator:uav_write
	wire          ch1_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                   // CH1_YN3_L_s1_translator_avalon_universal_slave_0_agent:m0_lock -> CH1_YN3_L_s1_translator:uav_lock
	wire          ch1_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_read;                                   // CH1_YN3_L_s1_translator_avalon_universal_slave_0_agent:m0_read -> CH1_YN3_L_s1_translator:uav_read
	wire   [31:0] ch1_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                               // CH1_YN3_L_s1_translator:uav_readdata -> CH1_YN3_L_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          ch1_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                          // CH1_YN3_L_s1_translator:uav_readdatavalid -> CH1_YN3_L_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          ch1_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                            // CH1_YN3_L_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> CH1_YN3_L_s1_translator:uav_debugaccess
	wire    [3:0] ch1_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                             // CH1_YN3_L_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> CH1_YN3_L_s1_translator:uav_byteenable
	wire          ch1_yn3_l_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                     // CH1_YN3_L_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> CH1_YN3_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          ch1_yn3_l_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                           // CH1_YN3_L_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> CH1_YN3_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          ch1_yn3_l_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                   // CH1_YN3_L_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> CH1_YN3_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] ch1_yn3_l_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                            // CH1_YN3_L_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> CH1_YN3_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          ch1_yn3_l_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                           // CH1_YN3_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> CH1_YN3_L_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          ch1_yn3_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                  // CH1_YN3_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> CH1_YN3_L_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          ch1_yn3_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                        // CH1_YN3_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> CH1_YN3_L_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          ch1_yn3_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                // CH1_YN3_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> CH1_YN3_L_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] ch1_yn3_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                         // CH1_YN3_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> CH1_YN3_L_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          ch1_yn3_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                        // CH1_YN3_L_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> CH1_YN3_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          ch1_yn3_l_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                      // CH1_YN3_L_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> CH1_YN3_L_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] ch1_yn3_l_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                       // CH1_YN3_L_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> CH1_YN3_L_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          ch1_yn3_l_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                      // CH1_YN3_L_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> CH1_YN3_L_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          ch2_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                        // CH2_TIMER_RST_s1_translator:uav_waitrequest -> CH2_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] ch2_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                         // CH2_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> CH2_TIMER_RST_s1_translator:uav_burstcount
	wire   [31:0] ch2_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                          // CH2_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> CH2_TIMER_RST_s1_translator:uav_writedata
	wire   [21:0] ch2_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_address;                            // CH2_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:m0_address -> CH2_TIMER_RST_s1_translator:uav_address
	wire          ch2_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_write;                              // CH2_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:m0_write -> CH2_TIMER_RST_s1_translator:uav_write
	wire          ch2_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_lock;                               // CH2_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:m0_lock -> CH2_TIMER_RST_s1_translator:uav_lock
	wire          ch2_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_read;                               // CH2_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:m0_read -> CH2_TIMER_RST_s1_translator:uav_read
	wire   [31:0] ch2_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                           // CH2_TIMER_RST_s1_translator:uav_readdata -> CH2_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          ch2_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                      // CH2_TIMER_RST_s1_translator:uav_readdatavalid -> CH2_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          ch2_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                        // CH2_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> CH2_TIMER_RST_s1_translator:uav_debugaccess
	wire    [3:0] ch2_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                         // CH2_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> CH2_TIMER_RST_s1_translator:uav_byteenable
	wire          ch2_timer_rst_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                 // CH2_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> CH2_TIMER_RST_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          ch2_timer_rst_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                       // CH2_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> CH2_TIMER_RST_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          ch2_timer_rst_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;               // CH2_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> CH2_TIMER_RST_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] ch2_timer_rst_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                        // CH2_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> CH2_TIMER_RST_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          ch2_timer_rst_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                       // CH2_TIMER_RST_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> CH2_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          ch2_timer_rst_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;              // CH2_TIMER_RST_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> CH2_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          ch2_timer_rst_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                    // CH2_TIMER_RST_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> CH2_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          ch2_timer_rst_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;            // CH2_TIMER_RST_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> CH2_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] ch2_timer_rst_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                     // CH2_TIMER_RST_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> CH2_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          ch2_timer_rst_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                    // CH2_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> CH2_TIMER_RST_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          ch2_timer_rst_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                  // CH2_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> CH2_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] ch2_timer_rst_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                   // CH2_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> CH2_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          ch2_timer_rst_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                  // CH2_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> CH2_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          ch2_thresh_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                           // CH2_THRESH_s1_translator:uav_waitrequest -> CH2_THRESH_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] ch2_thresh_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                            // CH2_THRESH_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> CH2_THRESH_s1_translator:uav_burstcount
	wire   [31:0] ch2_thresh_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                             // CH2_THRESH_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> CH2_THRESH_s1_translator:uav_writedata
	wire   [21:0] ch2_thresh_s1_translator_avalon_universal_slave_0_agent_m0_address;                               // CH2_THRESH_s1_translator_avalon_universal_slave_0_agent:m0_address -> CH2_THRESH_s1_translator:uav_address
	wire          ch2_thresh_s1_translator_avalon_universal_slave_0_agent_m0_write;                                 // CH2_THRESH_s1_translator_avalon_universal_slave_0_agent:m0_write -> CH2_THRESH_s1_translator:uav_write
	wire          ch2_thresh_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                  // CH2_THRESH_s1_translator_avalon_universal_slave_0_agent:m0_lock -> CH2_THRESH_s1_translator:uav_lock
	wire          ch2_thresh_s1_translator_avalon_universal_slave_0_agent_m0_read;                                  // CH2_THRESH_s1_translator_avalon_universal_slave_0_agent:m0_read -> CH2_THRESH_s1_translator:uav_read
	wire   [31:0] ch2_thresh_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                              // CH2_THRESH_s1_translator:uav_readdata -> CH2_THRESH_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          ch2_thresh_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                         // CH2_THRESH_s1_translator:uav_readdatavalid -> CH2_THRESH_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          ch2_thresh_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                           // CH2_THRESH_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> CH2_THRESH_s1_translator:uav_debugaccess
	wire    [3:0] ch2_thresh_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                            // CH2_THRESH_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> CH2_THRESH_s1_translator:uav_byteenable
	wire          ch2_thresh_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                    // CH2_THRESH_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> CH2_THRESH_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          ch2_thresh_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                          // CH2_THRESH_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> CH2_THRESH_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          ch2_thresh_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                  // CH2_THRESH_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> CH2_THRESH_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] ch2_thresh_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                           // CH2_THRESH_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> CH2_THRESH_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          ch2_thresh_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                          // CH2_THRESH_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> CH2_THRESH_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          ch2_thresh_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                 // CH2_THRESH_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> CH2_THRESH_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          ch2_thresh_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                       // CH2_THRESH_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> CH2_THRESH_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          ch2_thresh_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;               // CH2_THRESH_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> CH2_THRESH_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] ch2_thresh_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                        // CH2_THRESH_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> CH2_THRESH_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          ch2_thresh_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                       // CH2_THRESH_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> CH2_THRESH_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          ch2_thresh_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                     // CH2_THRESH_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> CH2_THRESH_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] ch2_thresh_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                      // CH2_THRESH_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> CH2_THRESH_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          ch2_thresh_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                     // CH2_THRESH_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> CH2_THRESH_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          ch2_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                          // CH2_RD_PEAK_s1_translator:uav_waitrequest -> CH2_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] ch2_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                           // CH2_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> CH2_RD_PEAK_s1_translator:uav_burstcount
	wire   [31:0] ch2_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                            // CH2_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> CH2_RD_PEAK_s1_translator:uav_writedata
	wire   [21:0] ch2_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_address;                              // CH2_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:m0_address -> CH2_RD_PEAK_s1_translator:uav_address
	wire          ch2_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_write;                                // CH2_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:m0_write -> CH2_RD_PEAK_s1_translator:uav_write
	wire          ch2_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                 // CH2_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:m0_lock -> CH2_RD_PEAK_s1_translator:uav_lock
	wire          ch2_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_read;                                 // CH2_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:m0_read -> CH2_RD_PEAK_s1_translator:uav_read
	wire   [31:0] ch2_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                             // CH2_RD_PEAK_s1_translator:uav_readdata -> CH2_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          ch2_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                        // CH2_RD_PEAK_s1_translator:uav_readdatavalid -> CH2_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          ch2_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                          // CH2_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> CH2_RD_PEAK_s1_translator:uav_debugaccess
	wire    [3:0] ch2_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                           // CH2_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> CH2_RD_PEAK_s1_translator:uav_byteenable
	wire          ch2_rd_peak_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                   // CH2_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> CH2_RD_PEAK_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          ch2_rd_peak_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                         // CH2_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> CH2_RD_PEAK_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          ch2_rd_peak_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                 // CH2_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> CH2_RD_PEAK_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] ch2_rd_peak_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                          // CH2_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> CH2_RD_PEAK_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          ch2_rd_peak_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                         // CH2_RD_PEAK_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> CH2_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          ch2_rd_peak_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                // CH2_RD_PEAK_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> CH2_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          ch2_rd_peak_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                      // CH2_RD_PEAK_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> CH2_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          ch2_rd_peak_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;              // CH2_RD_PEAK_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> CH2_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] ch2_rd_peak_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                       // CH2_RD_PEAK_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> CH2_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          ch2_rd_peak_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                      // CH2_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> CH2_RD_PEAK_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          ch2_rd_peak_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                    // CH2_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> CH2_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] ch2_rd_peak_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                     // CH2_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> CH2_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          ch2_rd_peak_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                    // CH2_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> CH2_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          ch2_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                       // CH2_PEAK_FOUND_s1_translator:uav_waitrequest -> CH2_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] ch2_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                        // CH2_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> CH2_PEAK_FOUND_s1_translator:uav_burstcount
	wire   [31:0] ch2_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                         // CH2_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> CH2_PEAK_FOUND_s1_translator:uav_writedata
	wire   [21:0] ch2_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_address;                           // CH2_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:m0_address -> CH2_PEAK_FOUND_s1_translator:uav_address
	wire          ch2_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_write;                             // CH2_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:m0_write -> CH2_PEAK_FOUND_s1_translator:uav_write
	wire          ch2_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_lock;                              // CH2_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:m0_lock -> CH2_PEAK_FOUND_s1_translator:uav_lock
	wire          ch2_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_read;                              // CH2_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:m0_read -> CH2_PEAK_FOUND_s1_translator:uav_read
	wire   [31:0] ch2_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                          // CH2_PEAK_FOUND_s1_translator:uav_readdata -> CH2_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          ch2_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                     // CH2_PEAK_FOUND_s1_translator:uav_readdatavalid -> CH2_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          ch2_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                       // CH2_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> CH2_PEAK_FOUND_s1_translator:uav_debugaccess
	wire    [3:0] ch2_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                        // CH2_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> CH2_PEAK_FOUND_s1_translator:uav_byteenable
	wire          ch2_peak_found_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                // CH2_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> CH2_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          ch2_peak_found_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                      // CH2_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> CH2_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          ch2_peak_found_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;              // CH2_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> CH2_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] ch2_peak_found_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                       // CH2_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> CH2_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          ch2_peak_found_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                      // CH2_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> CH2_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          ch2_peak_found_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;             // CH2_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> CH2_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          ch2_peak_found_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                   // CH2_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> CH2_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          ch2_peak_found_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;           // CH2_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> CH2_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] ch2_peak_found_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                    // CH2_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> CH2_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          ch2_peak_found_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                   // CH2_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> CH2_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          ch2_peak_found_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                 // CH2_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> CH2_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] ch2_peak_found_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                  // CH2_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> CH2_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          ch2_peak_found_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                 // CH2_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> CH2_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          ch2_time_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                             // CH2_TIME_s1_translator:uav_waitrequest -> CH2_TIME_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] ch2_time_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                              // CH2_TIME_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> CH2_TIME_s1_translator:uav_burstcount
	wire   [31:0] ch2_time_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                               // CH2_TIME_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> CH2_TIME_s1_translator:uav_writedata
	wire   [21:0] ch2_time_s1_translator_avalon_universal_slave_0_agent_m0_address;                                 // CH2_TIME_s1_translator_avalon_universal_slave_0_agent:m0_address -> CH2_TIME_s1_translator:uav_address
	wire          ch2_time_s1_translator_avalon_universal_slave_0_agent_m0_write;                                   // CH2_TIME_s1_translator_avalon_universal_slave_0_agent:m0_write -> CH2_TIME_s1_translator:uav_write
	wire          ch2_time_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                    // CH2_TIME_s1_translator_avalon_universal_slave_0_agent:m0_lock -> CH2_TIME_s1_translator:uav_lock
	wire          ch2_time_s1_translator_avalon_universal_slave_0_agent_m0_read;                                    // CH2_TIME_s1_translator_avalon_universal_slave_0_agent:m0_read -> CH2_TIME_s1_translator:uav_read
	wire   [31:0] ch2_time_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                // CH2_TIME_s1_translator:uav_readdata -> CH2_TIME_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          ch2_time_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                           // CH2_TIME_s1_translator:uav_readdatavalid -> CH2_TIME_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          ch2_time_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                             // CH2_TIME_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> CH2_TIME_s1_translator:uav_debugaccess
	wire    [3:0] ch2_time_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                              // CH2_TIME_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> CH2_TIME_s1_translator:uav_byteenable
	wire          ch2_time_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                      // CH2_TIME_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> CH2_TIME_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          ch2_time_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                            // CH2_TIME_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> CH2_TIME_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          ch2_time_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                    // CH2_TIME_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> CH2_TIME_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] ch2_time_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                             // CH2_TIME_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> CH2_TIME_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          ch2_time_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                            // CH2_TIME_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> CH2_TIME_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          ch2_time_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                   // CH2_TIME_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> CH2_TIME_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          ch2_time_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                         // CH2_TIME_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> CH2_TIME_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          ch2_time_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                 // CH2_TIME_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> CH2_TIME_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] ch2_time_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                          // CH2_TIME_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> CH2_TIME_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          ch2_time_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                         // CH2_TIME_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> CH2_TIME_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          ch2_time_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                       // CH2_TIME_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> CH2_TIME_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] ch2_time_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                        // CH2_TIME_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> CH2_TIME_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          ch2_time_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                       // CH2_TIME_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> CH2_TIME_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          ch2_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                            // CH2_YN1_U_s1_translator:uav_waitrequest -> CH2_YN1_U_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] ch2_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                             // CH2_YN1_U_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> CH2_YN1_U_s1_translator:uav_burstcount
	wire   [31:0] ch2_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                              // CH2_YN1_U_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> CH2_YN1_U_s1_translator:uav_writedata
	wire   [21:0] ch2_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_address;                                // CH2_YN1_U_s1_translator_avalon_universal_slave_0_agent:m0_address -> CH2_YN1_U_s1_translator:uav_address
	wire          ch2_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_write;                                  // CH2_YN1_U_s1_translator_avalon_universal_slave_0_agent:m0_write -> CH2_YN1_U_s1_translator:uav_write
	wire          ch2_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                   // CH2_YN1_U_s1_translator_avalon_universal_slave_0_agent:m0_lock -> CH2_YN1_U_s1_translator:uav_lock
	wire          ch2_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_read;                                   // CH2_YN1_U_s1_translator_avalon_universal_slave_0_agent:m0_read -> CH2_YN1_U_s1_translator:uav_read
	wire   [31:0] ch2_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                               // CH2_YN1_U_s1_translator:uav_readdata -> CH2_YN1_U_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          ch2_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                          // CH2_YN1_U_s1_translator:uav_readdatavalid -> CH2_YN1_U_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          ch2_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                            // CH2_YN1_U_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> CH2_YN1_U_s1_translator:uav_debugaccess
	wire    [3:0] ch2_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                             // CH2_YN1_U_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> CH2_YN1_U_s1_translator:uav_byteenable
	wire          ch2_yn1_u_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                     // CH2_YN1_U_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> CH2_YN1_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          ch2_yn1_u_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                           // CH2_YN1_U_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> CH2_YN1_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          ch2_yn1_u_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                   // CH2_YN1_U_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> CH2_YN1_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] ch2_yn1_u_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                            // CH2_YN1_U_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> CH2_YN1_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          ch2_yn1_u_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                           // CH2_YN1_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> CH2_YN1_U_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          ch2_yn1_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                  // CH2_YN1_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> CH2_YN1_U_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          ch2_yn1_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                        // CH2_YN1_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> CH2_YN1_U_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          ch2_yn1_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                // CH2_YN1_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> CH2_YN1_U_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] ch2_yn1_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                         // CH2_YN1_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> CH2_YN1_U_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          ch2_yn1_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                        // CH2_YN1_U_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> CH2_YN1_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          ch2_yn1_u_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                      // CH2_YN1_U_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> CH2_YN1_U_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] ch2_yn1_u_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                       // CH2_YN1_U_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> CH2_YN1_U_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          ch2_yn1_u_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                      // CH2_YN1_U_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> CH2_YN1_U_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          ch2_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                           // CH2_YN1_MU_s1_translator:uav_waitrequest -> CH2_YN1_MU_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] ch2_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                            // CH2_YN1_MU_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> CH2_YN1_MU_s1_translator:uav_burstcount
	wire   [31:0] ch2_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                             // CH2_YN1_MU_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> CH2_YN1_MU_s1_translator:uav_writedata
	wire   [21:0] ch2_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_address;                               // CH2_YN1_MU_s1_translator_avalon_universal_slave_0_agent:m0_address -> CH2_YN1_MU_s1_translator:uav_address
	wire          ch2_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_write;                                 // CH2_YN1_MU_s1_translator_avalon_universal_slave_0_agent:m0_write -> CH2_YN1_MU_s1_translator:uav_write
	wire          ch2_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                  // CH2_YN1_MU_s1_translator_avalon_universal_slave_0_agent:m0_lock -> CH2_YN1_MU_s1_translator:uav_lock
	wire          ch2_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_read;                                  // CH2_YN1_MU_s1_translator_avalon_universal_slave_0_agent:m0_read -> CH2_YN1_MU_s1_translator:uav_read
	wire   [31:0] ch2_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                              // CH2_YN1_MU_s1_translator:uav_readdata -> CH2_YN1_MU_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          ch2_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                         // CH2_YN1_MU_s1_translator:uav_readdatavalid -> CH2_YN1_MU_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          ch2_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                           // CH2_YN1_MU_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> CH2_YN1_MU_s1_translator:uav_debugaccess
	wire    [3:0] ch2_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                            // CH2_YN1_MU_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> CH2_YN1_MU_s1_translator:uav_byteenable
	wire          ch2_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                    // CH2_YN1_MU_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> CH2_YN1_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          ch2_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                          // CH2_YN1_MU_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> CH2_YN1_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          ch2_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                  // CH2_YN1_MU_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> CH2_YN1_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] ch2_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                           // CH2_YN1_MU_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> CH2_YN1_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          ch2_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                          // CH2_YN1_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> CH2_YN1_MU_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          ch2_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                 // CH2_YN1_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> CH2_YN1_MU_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          ch2_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                       // CH2_YN1_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> CH2_YN1_MU_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          ch2_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;               // CH2_YN1_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> CH2_YN1_MU_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] ch2_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                        // CH2_YN1_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> CH2_YN1_MU_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          ch2_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                       // CH2_YN1_MU_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> CH2_YN1_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          ch2_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                     // CH2_YN1_MU_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> CH2_YN1_MU_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] ch2_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                      // CH2_YN1_MU_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> CH2_YN1_MU_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          ch2_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                     // CH2_YN1_MU_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> CH2_YN1_MU_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          ch2_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                           // CH2_YN1_ML_s1_translator:uav_waitrequest -> CH2_YN1_ML_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] ch2_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                            // CH2_YN1_ML_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> CH2_YN1_ML_s1_translator:uav_burstcount
	wire   [31:0] ch2_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                             // CH2_YN1_ML_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> CH2_YN1_ML_s1_translator:uav_writedata
	wire   [21:0] ch2_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_address;                               // CH2_YN1_ML_s1_translator_avalon_universal_slave_0_agent:m0_address -> CH2_YN1_ML_s1_translator:uav_address
	wire          ch2_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_write;                                 // CH2_YN1_ML_s1_translator_avalon_universal_slave_0_agent:m0_write -> CH2_YN1_ML_s1_translator:uav_write
	wire          ch2_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                  // CH2_YN1_ML_s1_translator_avalon_universal_slave_0_agent:m0_lock -> CH2_YN1_ML_s1_translator:uav_lock
	wire          ch2_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_read;                                  // CH2_YN1_ML_s1_translator_avalon_universal_slave_0_agent:m0_read -> CH2_YN1_ML_s1_translator:uav_read
	wire   [31:0] ch2_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                              // CH2_YN1_ML_s1_translator:uav_readdata -> CH2_YN1_ML_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          ch2_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                         // CH2_YN1_ML_s1_translator:uav_readdatavalid -> CH2_YN1_ML_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          ch2_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                           // CH2_YN1_ML_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> CH2_YN1_ML_s1_translator:uav_debugaccess
	wire    [3:0] ch2_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                            // CH2_YN1_ML_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> CH2_YN1_ML_s1_translator:uav_byteenable
	wire          ch2_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                    // CH2_YN1_ML_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> CH2_YN1_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          ch2_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                          // CH2_YN1_ML_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> CH2_YN1_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          ch2_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                  // CH2_YN1_ML_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> CH2_YN1_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] ch2_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                           // CH2_YN1_ML_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> CH2_YN1_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          ch2_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                          // CH2_YN1_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> CH2_YN1_ML_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          ch2_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                 // CH2_YN1_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> CH2_YN1_ML_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          ch2_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                       // CH2_YN1_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> CH2_YN1_ML_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          ch2_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;               // CH2_YN1_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> CH2_YN1_ML_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] ch2_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                        // CH2_YN1_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> CH2_YN1_ML_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          ch2_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                       // CH2_YN1_ML_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> CH2_YN1_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          ch2_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                     // CH2_YN1_ML_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> CH2_YN1_ML_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] ch2_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                      // CH2_YN1_ML_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> CH2_YN1_ML_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          ch2_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                     // CH2_YN1_ML_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> CH2_YN1_ML_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          ch2_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                            // CH2_YN1_L_s1_translator:uav_waitrequest -> CH2_YN1_L_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] ch2_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                             // CH2_YN1_L_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> CH2_YN1_L_s1_translator:uav_burstcount
	wire   [31:0] ch2_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                              // CH2_YN1_L_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> CH2_YN1_L_s1_translator:uav_writedata
	wire   [21:0] ch2_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_address;                                // CH2_YN1_L_s1_translator_avalon_universal_slave_0_agent:m0_address -> CH2_YN1_L_s1_translator:uav_address
	wire          ch2_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_write;                                  // CH2_YN1_L_s1_translator_avalon_universal_slave_0_agent:m0_write -> CH2_YN1_L_s1_translator:uav_write
	wire          ch2_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                   // CH2_YN1_L_s1_translator_avalon_universal_slave_0_agent:m0_lock -> CH2_YN1_L_s1_translator:uav_lock
	wire          ch2_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_read;                                   // CH2_YN1_L_s1_translator_avalon_universal_slave_0_agent:m0_read -> CH2_YN1_L_s1_translator:uav_read
	wire   [31:0] ch2_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                               // CH2_YN1_L_s1_translator:uav_readdata -> CH2_YN1_L_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          ch2_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                          // CH2_YN1_L_s1_translator:uav_readdatavalid -> CH2_YN1_L_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          ch2_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                            // CH2_YN1_L_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> CH2_YN1_L_s1_translator:uav_debugaccess
	wire    [3:0] ch2_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                             // CH2_YN1_L_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> CH2_YN1_L_s1_translator:uav_byteenable
	wire          ch2_yn1_l_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                     // CH2_YN1_L_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> CH2_YN1_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          ch2_yn1_l_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                           // CH2_YN1_L_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> CH2_YN1_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          ch2_yn1_l_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                   // CH2_YN1_L_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> CH2_YN1_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] ch2_yn1_l_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                            // CH2_YN1_L_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> CH2_YN1_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          ch2_yn1_l_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                           // CH2_YN1_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> CH2_YN1_L_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          ch2_yn1_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                  // CH2_YN1_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> CH2_YN1_L_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          ch2_yn1_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                        // CH2_YN1_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> CH2_YN1_L_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          ch2_yn1_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                // CH2_YN1_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> CH2_YN1_L_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] ch2_yn1_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                         // CH2_YN1_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> CH2_YN1_L_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          ch2_yn1_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                        // CH2_YN1_L_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> CH2_YN1_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          ch2_yn1_l_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                      // CH2_YN1_L_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> CH2_YN1_L_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] ch2_yn1_l_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                       // CH2_YN1_L_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> CH2_YN1_L_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          ch2_yn1_l_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                      // CH2_YN1_L_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> CH2_YN1_L_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          ch2_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                            // CH2_YN2_U_s1_translator:uav_waitrequest -> CH2_YN2_U_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] ch2_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                             // CH2_YN2_U_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> CH2_YN2_U_s1_translator:uav_burstcount
	wire   [31:0] ch2_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                              // CH2_YN2_U_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> CH2_YN2_U_s1_translator:uav_writedata
	wire   [21:0] ch2_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_address;                                // CH2_YN2_U_s1_translator_avalon_universal_slave_0_agent:m0_address -> CH2_YN2_U_s1_translator:uav_address
	wire          ch2_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_write;                                  // CH2_YN2_U_s1_translator_avalon_universal_slave_0_agent:m0_write -> CH2_YN2_U_s1_translator:uav_write
	wire          ch2_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                   // CH2_YN2_U_s1_translator_avalon_universal_slave_0_agent:m0_lock -> CH2_YN2_U_s1_translator:uav_lock
	wire          ch2_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_read;                                   // CH2_YN2_U_s1_translator_avalon_universal_slave_0_agent:m0_read -> CH2_YN2_U_s1_translator:uav_read
	wire   [31:0] ch2_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                               // CH2_YN2_U_s1_translator:uav_readdata -> CH2_YN2_U_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          ch2_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                          // CH2_YN2_U_s1_translator:uav_readdatavalid -> CH2_YN2_U_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          ch2_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                            // CH2_YN2_U_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> CH2_YN2_U_s1_translator:uav_debugaccess
	wire    [3:0] ch2_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                             // CH2_YN2_U_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> CH2_YN2_U_s1_translator:uav_byteenable
	wire          ch2_yn2_u_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                     // CH2_YN2_U_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> CH2_YN2_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          ch2_yn2_u_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                           // CH2_YN2_U_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> CH2_YN2_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          ch2_yn2_u_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                   // CH2_YN2_U_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> CH2_YN2_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] ch2_yn2_u_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                            // CH2_YN2_U_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> CH2_YN2_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          ch2_yn2_u_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                           // CH2_YN2_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> CH2_YN2_U_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          ch2_yn2_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                  // CH2_YN2_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> CH2_YN2_U_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          ch2_yn2_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                        // CH2_YN2_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> CH2_YN2_U_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          ch2_yn2_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                // CH2_YN2_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> CH2_YN2_U_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] ch2_yn2_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                         // CH2_YN2_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> CH2_YN2_U_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          ch2_yn2_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                        // CH2_YN2_U_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> CH2_YN2_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          ch2_yn2_u_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                      // CH2_YN2_U_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> CH2_YN2_U_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] ch2_yn2_u_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                       // CH2_YN2_U_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> CH2_YN2_U_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          ch2_yn2_u_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                      // CH2_YN2_U_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> CH2_YN2_U_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          ch2_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                           // CH2_YN2_MU_s1_translator:uav_waitrequest -> CH2_YN2_MU_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] ch2_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                            // CH2_YN2_MU_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> CH2_YN2_MU_s1_translator:uav_burstcount
	wire   [31:0] ch2_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                             // CH2_YN2_MU_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> CH2_YN2_MU_s1_translator:uav_writedata
	wire   [21:0] ch2_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_address;                               // CH2_YN2_MU_s1_translator_avalon_universal_slave_0_agent:m0_address -> CH2_YN2_MU_s1_translator:uav_address
	wire          ch2_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_write;                                 // CH2_YN2_MU_s1_translator_avalon_universal_slave_0_agent:m0_write -> CH2_YN2_MU_s1_translator:uav_write
	wire          ch2_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                  // CH2_YN2_MU_s1_translator_avalon_universal_slave_0_agent:m0_lock -> CH2_YN2_MU_s1_translator:uav_lock
	wire          ch2_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_read;                                  // CH2_YN2_MU_s1_translator_avalon_universal_slave_0_agent:m0_read -> CH2_YN2_MU_s1_translator:uav_read
	wire   [31:0] ch2_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                              // CH2_YN2_MU_s1_translator:uav_readdata -> CH2_YN2_MU_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          ch2_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                         // CH2_YN2_MU_s1_translator:uav_readdatavalid -> CH2_YN2_MU_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          ch2_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                           // CH2_YN2_MU_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> CH2_YN2_MU_s1_translator:uav_debugaccess
	wire    [3:0] ch2_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                            // CH2_YN2_MU_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> CH2_YN2_MU_s1_translator:uav_byteenable
	wire          ch2_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                    // CH2_YN2_MU_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> CH2_YN2_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          ch2_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                          // CH2_YN2_MU_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> CH2_YN2_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          ch2_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                  // CH2_YN2_MU_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> CH2_YN2_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] ch2_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                           // CH2_YN2_MU_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> CH2_YN2_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          ch2_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                          // CH2_YN2_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> CH2_YN2_MU_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          ch2_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                 // CH2_YN2_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> CH2_YN2_MU_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          ch2_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                       // CH2_YN2_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> CH2_YN2_MU_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          ch2_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;               // CH2_YN2_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> CH2_YN2_MU_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] ch2_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                        // CH2_YN2_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> CH2_YN2_MU_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          ch2_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                       // CH2_YN2_MU_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> CH2_YN2_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          ch2_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                     // CH2_YN2_MU_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> CH2_YN2_MU_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] ch2_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                      // CH2_YN2_MU_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> CH2_YN2_MU_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          ch2_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                     // CH2_YN2_MU_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> CH2_YN2_MU_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          ch2_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                           // CH2_YN2_ML_s1_translator:uav_waitrequest -> CH2_YN2_ML_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] ch2_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                            // CH2_YN2_ML_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> CH2_YN2_ML_s1_translator:uav_burstcount
	wire   [31:0] ch2_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                             // CH2_YN2_ML_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> CH2_YN2_ML_s1_translator:uav_writedata
	wire   [21:0] ch2_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_address;                               // CH2_YN2_ML_s1_translator_avalon_universal_slave_0_agent:m0_address -> CH2_YN2_ML_s1_translator:uav_address
	wire          ch2_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_write;                                 // CH2_YN2_ML_s1_translator_avalon_universal_slave_0_agent:m0_write -> CH2_YN2_ML_s1_translator:uav_write
	wire          ch2_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                  // CH2_YN2_ML_s1_translator_avalon_universal_slave_0_agent:m0_lock -> CH2_YN2_ML_s1_translator:uav_lock
	wire          ch2_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_read;                                  // CH2_YN2_ML_s1_translator_avalon_universal_slave_0_agent:m0_read -> CH2_YN2_ML_s1_translator:uav_read
	wire   [31:0] ch2_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                              // CH2_YN2_ML_s1_translator:uav_readdata -> CH2_YN2_ML_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          ch2_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                         // CH2_YN2_ML_s1_translator:uav_readdatavalid -> CH2_YN2_ML_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          ch2_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                           // CH2_YN2_ML_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> CH2_YN2_ML_s1_translator:uav_debugaccess
	wire    [3:0] ch2_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                            // CH2_YN2_ML_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> CH2_YN2_ML_s1_translator:uav_byteenable
	wire          ch2_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                    // CH2_YN2_ML_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> CH2_YN2_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          ch2_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                          // CH2_YN2_ML_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> CH2_YN2_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          ch2_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                  // CH2_YN2_ML_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> CH2_YN2_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] ch2_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                           // CH2_YN2_ML_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> CH2_YN2_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          ch2_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                          // CH2_YN2_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> CH2_YN2_ML_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          ch2_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                 // CH2_YN2_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> CH2_YN2_ML_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          ch2_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                       // CH2_YN2_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> CH2_YN2_ML_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          ch2_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;               // CH2_YN2_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> CH2_YN2_ML_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] ch2_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                        // CH2_YN2_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> CH2_YN2_ML_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          ch2_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                       // CH2_YN2_ML_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> CH2_YN2_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          ch2_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                     // CH2_YN2_ML_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> CH2_YN2_ML_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] ch2_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                      // CH2_YN2_ML_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> CH2_YN2_ML_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          ch2_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                     // CH2_YN2_ML_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> CH2_YN2_ML_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          ch2_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                            // CH2_YN2_L_s1_translator:uav_waitrequest -> CH2_YN2_L_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] ch2_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                             // CH2_YN2_L_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> CH2_YN2_L_s1_translator:uav_burstcount
	wire   [31:0] ch2_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                              // CH2_YN2_L_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> CH2_YN2_L_s1_translator:uav_writedata
	wire   [21:0] ch2_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_address;                                // CH2_YN2_L_s1_translator_avalon_universal_slave_0_agent:m0_address -> CH2_YN2_L_s1_translator:uav_address
	wire          ch2_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_write;                                  // CH2_YN2_L_s1_translator_avalon_universal_slave_0_agent:m0_write -> CH2_YN2_L_s1_translator:uav_write
	wire          ch2_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                   // CH2_YN2_L_s1_translator_avalon_universal_slave_0_agent:m0_lock -> CH2_YN2_L_s1_translator:uav_lock
	wire          ch2_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_read;                                   // CH2_YN2_L_s1_translator_avalon_universal_slave_0_agent:m0_read -> CH2_YN2_L_s1_translator:uav_read
	wire   [31:0] ch2_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                               // CH2_YN2_L_s1_translator:uav_readdata -> CH2_YN2_L_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          ch2_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                          // CH2_YN2_L_s1_translator:uav_readdatavalid -> CH2_YN2_L_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          ch2_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                            // CH2_YN2_L_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> CH2_YN2_L_s1_translator:uav_debugaccess
	wire    [3:0] ch2_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                             // CH2_YN2_L_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> CH2_YN2_L_s1_translator:uav_byteenable
	wire          ch2_yn2_l_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                     // CH2_YN2_L_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> CH2_YN2_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          ch2_yn2_l_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                           // CH2_YN2_L_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> CH2_YN2_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          ch2_yn2_l_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                   // CH2_YN2_L_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> CH2_YN2_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] ch2_yn2_l_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                            // CH2_YN2_L_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> CH2_YN2_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          ch2_yn2_l_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                           // CH2_YN2_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> CH2_YN2_L_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          ch2_yn2_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                  // CH2_YN2_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> CH2_YN2_L_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          ch2_yn2_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                        // CH2_YN2_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> CH2_YN2_L_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          ch2_yn2_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                // CH2_YN2_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> CH2_YN2_L_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] ch2_yn2_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                         // CH2_YN2_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> CH2_YN2_L_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          ch2_yn2_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                        // CH2_YN2_L_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> CH2_YN2_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          ch2_yn2_l_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                      // CH2_YN2_L_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> CH2_YN2_L_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] ch2_yn2_l_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                       // CH2_YN2_L_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> CH2_YN2_L_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          ch2_yn2_l_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                      // CH2_YN2_L_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> CH2_YN2_L_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          ch2_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                            // CH2_YN3_U_s1_translator:uav_waitrequest -> CH2_YN3_U_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] ch2_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                             // CH2_YN3_U_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> CH2_YN3_U_s1_translator:uav_burstcount
	wire   [31:0] ch2_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                              // CH2_YN3_U_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> CH2_YN3_U_s1_translator:uav_writedata
	wire   [21:0] ch2_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_address;                                // CH2_YN3_U_s1_translator_avalon_universal_slave_0_agent:m0_address -> CH2_YN3_U_s1_translator:uav_address
	wire          ch2_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_write;                                  // CH2_YN3_U_s1_translator_avalon_universal_slave_0_agent:m0_write -> CH2_YN3_U_s1_translator:uav_write
	wire          ch2_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                   // CH2_YN3_U_s1_translator_avalon_universal_slave_0_agent:m0_lock -> CH2_YN3_U_s1_translator:uav_lock
	wire          ch2_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_read;                                   // CH2_YN3_U_s1_translator_avalon_universal_slave_0_agent:m0_read -> CH2_YN3_U_s1_translator:uav_read
	wire   [31:0] ch2_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                               // CH2_YN3_U_s1_translator:uav_readdata -> CH2_YN3_U_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          ch2_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                          // CH2_YN3_U_s1_translator:uav_readdatavalid -> CH2_YN3_U_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          ch2_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                            // CH2_YN3_U_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> CH2_YN3_U_s1_translator:uav_debugaccess
	wire    [3:0] ch2_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                             // CH2_YN3_U_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> CH2_YN3_U_s1_translator:uav_byteenable
	wire          ch2_yn3_u_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                     // CH2_YN3_U_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> CH2_YN3_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          ch2_yn3_u_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                           // CH2_YN3_U_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> CH2_YN3_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          ch2_yn3_u_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                   // CH2_YN3_U_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> CH2_YN3_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] ch2_yn3_u_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                            // CH2_YN3_U_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> CH2_YN3_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          ch2_yn3_u_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                           // CH2_YN3_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> CH2_YN3_U_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          ch2_yn3_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                  // CH2_YN3_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> CH2_YN3_U_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          ch2_yn3_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                        // CH2_YN3_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> CH2_YN3_U_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          ch2_yn3_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                // CH2_YN3_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> CH2_YN3_U_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] ch2_yn3_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                         // CH2_YN3_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> CH2_YN3_U_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          ch2_yn3_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                        // CH2_YN3_U_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> CH2_YN3_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          ch2_yn3_u_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                      // CH2_YN3_U_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> CH2_YN3_U_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] ch2_yn3_u_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                       // CH2_YN3_U_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> CH2_YN3_U_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          ch2_yn3_u_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                      // CH2_YN3_U_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> CH2_YN3_U_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          ch2_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                           // CH2_YN3_MU_s1_translator:uav_waitrequest -> CH2_YN3_MU_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] ch2_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                            // CH2_YN3_MU_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> CH2_YN3_MU_s1_translator:uav_burstcount
	wire   [31:0] ch2_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                             // CH2_YN3_MU_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> CH2_YN3_MU_s1_translator:uav_writedata
	wire   [21:0] ch2_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_address;                               // CH2_YN3_MU_s1_translator_avalon_universal_slave_0_agent:m0_address -> CH2_YN3_MU_s1_translator:uav_address
	wire          ch2_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_write;                                 // CH2_YN3_MU_s1_translator_avalon_universal_slave_0_agent:m0_write -> CH2_YN3_MU_s1_translator:uav_write
	wire          ch2_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                  // CH2_YN3_MU_s1_translator_avalon_universal_slave_0_agent:m0_lock -> CH2_YN3_MU_s1_translator:uav_lock
	wire          ch2_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_read;                                  // CH2_YN3_MU_s1_translator_avalon_universal_slave_0_agent:m0_read -> CH2_YN3_MU_s1_translator:uav_read
	wire   [31:0] ch2_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                              // CH2_YN3_MU_s1_translator:uav_readdata -> CH2_YN3_MU_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          ch2_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                         // CH2_YN3_MU_s1_translator:uav_readdatavalid -> CH2_YN3_MU_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          ch2_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                           // CH2_YN3_MU_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> CH2_YN3_MU_s1_translator:uav_debugaccess
	wire    [3:0] ch2_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                            // CH2_YN3_MU_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> CH2_YN3_MU_s1_translator:uav_byteenable
	wire          ch2_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                    // CH2_YN3_MU_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> CH2_YN3_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          ch2_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                          // CH2_YN3_MU_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> CH2_YN3_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          ch2_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                  // CH2_YN3_MU_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> CH2_YN3_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] ch2_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                           // CH2_YN3_MU_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> CH2_YN3_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          ch2_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                          // CH2_YN3_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> CH2_YN3_MU_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          ch2_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                 // CH2_YN3_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> CH2_YN3_MU_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          ch2_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                       // CH2_YN3_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> CH2_YN3_MU_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          ch2_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;               // CH2_YN3_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> CH2_YN3_MU_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] ch2_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                        // CH2_YN3_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> CH2_YN3_MU_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          ch2_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                       // CH2_YN3_MU_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> CH2_YN3_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          ch2_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                     // CH2_YN3_MU_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> CH2_YN3_MU_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] ch2_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                      // CH2_YN3_MU_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> CH2_YN3_MU_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          ch2_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                     // CH2_YN3_MU_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> CH2_YN3_MU_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          ch2_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                           // CH2_YN3_ML_s1_translator:uav_waitrequest -> CH2_YN3_ML_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] ch2_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                            // CH2_YN3_ML_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> CH2_YN3_ML_s1_translator:uav_burstcount
	wire   [31:0] ch2_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                             // CH2_YN3_ML_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> CH2_YN3_ML_s1_translator:uav_writedata
	wire   [21:0] ch2_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_address;                               // CH2_YN3_ML_s1_translator_avalon_universal_slave_0_agent:m0_address -> CH2_YN3_ML_s1_translator:uav_address
	wire          ch2_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_write;                                 // CH2_YN3_ML_s1_translator_avalon_universal_slave_0_agent:m0_write -> CH2_YN3_ML_s1_translator:uav_write
	wire          ch2_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                  // CH2_YN3_ML_s1_translator_avalon_universal_slave_0_agent:m0_lock -> CH2_YN3_ML_s1_translator:uav_lock
	wire          ch2_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_read;                                  // CH2_YN3_ML_s1_translator_avalon_universal_slave_0_agent:m0_read -> CH2_YN3_ML_s1_translator:uav_read
	wire   [31:0] ch2_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                              // CH2_YN3_ML_s1_translator:uav_readdata -> CH2_YN3_ML_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          ch2_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                         // CH2_YN3_ML_s1_translator:uav_readdatavalid -> CH2_YN3_ML_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          ch2_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                           // CH2_YN3_ML_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> CH2_YN3_ML_s1_translator:uav_debugaccess
	wire    [3:0] ch2_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                            // CH2_YN3_ML_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> CH2_YN3_ML_s1_translator:uav_byteenable
	wire          ch2_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                    // CH2_YN3_ML_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> CH2_YN3_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          ch2_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                          // CH2_YN3_ML_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> CH2_YN3_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          ch2_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                  // CH2_YN3_ML_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> CH2_YN3_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] ch2_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                           // CH2_YN3_ML_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> CH2_YN3_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          ch2_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                          // CH2_YN3_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> CH2_YN3_ML_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          ch2_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                 // CH2_YN3_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> CH2_YN3_ML_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          ch2_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                       // CH2_YN3_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> CH2_YN3_ML_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          ch2_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;               // CH2_YN3_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> CH2_YN3_ML_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] ch2_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                        // CH2_YN3_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> CH2_YN3_ML_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          ch2_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                       // CH2_YN3_ML_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> CH2_YN3_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          ch2_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                     // CH2_YN3_ML_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> CH2_YN3_ML_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] ch2_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                      // CH2_YN3_ML_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> CH2_YN3_ML_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          ch2_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                     // CH2_YN3_ML_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> CH2_YN3_ML_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          ch2_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                            // CH2_YN3_L_s1_translator:uav_waitrequest -> CH2_YN3_L_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] ch2_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                             // CH2_YN3_L_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> CH2_YN3_L_s1_translator:uav_burstcount
	wire   [31:0] ch2_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                              // CH2_YN3_L_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> CH2_YN3_L_s1_translator:uav_writedata
	wire   [21:0] ch2_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_address;                                // CH2_YN3_L_s1_translator_avalon_universal_slave_0_agent:m0_address -> CH2_YN3_L_s1_translator:uav_address
	wire          ch2_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_write;                                  // CH2_YN3_L_s1_translator_avalon_universal_slave_0_agent:m0_write -> CH2_YN3_L_s1_translator:uav_write
	wire          ch2_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                   // CH2_YN3_L_s1_translator_avalon_universal_slave_0_agent:m0_lock -> CH2_YN3_L_s1_translator:uav_lock
	wire          ch2_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_read;                                   // CH2_YN3_L_s1_translator_avalon_universal_slave_0_agent:m0_read -> CH2_YN3_L_s1_translator:uav_read
	wire   [31:0] ch2_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                               // CH2_YN3_L_s1_translator:uav_readdata -> CH2_YN3_L_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          ch2_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                          // CH2_YN3_L_s1_translator:uav_readdatavalid -> CH2_YN3_L_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          ch2_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                            // CH2_YN3_L_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> CH2_YN3_L_s1_translator:uav_debugaccess
	wire    [3:0] ch2_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                             // CH2_YN3_L_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> CH2_YN3_L_s1_translator:uav_byteenable
	wire          ch2_yn3_l_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                     // CH2_YN3_L_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> CH2_YN3_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          ch2_yn3_l_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                           // CH2_YN3_L_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> CH2_YN3_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          ch2_yn3_l_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                   // CH2_YN3_L_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> CH2_YN3_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] ch2_yn3_l_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                            // CH2_YN3_L_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> CH2_YN3_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          ch2_yn3_l_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                           // CH2_YN3_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> CH2_YN3_L_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          ch2_yn3_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                  // CH2_YN3_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> CH2_YN3_L_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          ch2_yn3_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                        // CH2_YN3_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> CH2_YN3_L_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          ch2_yn3_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                // CH2_YN3_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> CH2_YN3_L_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] ch2_yn3_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                         // CH2_YN3_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> CH2_YN3_L_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          ch2_yn3_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                        // CH2_YN3_L_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> CH2_YN3_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          ch2_yn3_l_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                      // CH2_YN3_L_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> CH2_YN3_L_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] ch2_yn3_l_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                       // CH2_YN3_L_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> CH2_YN3_L_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          ch2_yn3_l_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                      // CH2_YN3_L_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> CH2_YN3_L_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          ch3_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                        // CH3_TIMER_RST_s1_translator:uav_waitrequest -> CH3_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] ch3_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                         // CH3_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> CH3_TIMER_RST_s1_translator:uav_burstcount
	wire   [31:0] ch3_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                          // CH3_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> CH3_TIMER_RST_s1_translator:uav_writedata
	wire   [21:0] ch3_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_address;                            // CH3_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:m0_address -> CH3_TIMER_RST_s1_translator:uav_address
	wire          ch3_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_write;                              // CH3_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:m0_write -> CH3_TIMER_RST_s1_translator:uav_write
	wire          ch3_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_lock;                               // CH3_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:m0_lock -> CH3_TIMER_RST_s1_translator:uav_lock
	wire          ch3_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_read;                               // CH3_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:m0_read -> CH3_TIMER_RST_s1_translator:uav_read
	wire   [31:0] ch3_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                           // CH3_TIMER_RST_s1_translator:uav_readdata -> CH3_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          ch3_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                      // CH3_TIMER_RST_s1_translator:uav_readdatavalid -> CH3_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          ch3_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                        // CH3_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> CH3_TIMER_RST_s1_translator:uav_debugaccess
	wire    [3:0] ch3_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                         // CH3_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> CH3_TIMER_RST_s1_translator:uav_byteenable
	wire          ch3_timer_rst_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                 // CH3_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> CH3_TIMER_RST_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          ch3_timer_rst_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                       // CH3_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> CH3_TIMER_RST_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          ch3_timer_rst_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;               // CH3_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> CH3_TIMER_RST_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] ch3_timer_rst_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                        // CH3_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> CH3_TIMER_RST_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          ch3_timer_rst_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                       // CH3_TIMER_RST_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> CH3_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          ch3_timer_rst_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;              // CH3_TIMER_RST_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> CH3_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          ch3_timer_rst_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                    // CH3_TIMER_RST_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> CH3_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          ch3_timer_rst_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;            // CH3_TIMER_RST_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> CH3_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] ch3_timer_rst_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                     // CH3_TIMER_RST_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> CH3_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          ch3_timer_rst_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                    // CH3_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> CH3_TIMER_RST_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          ch3_timer_rst_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                  // CH3_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> CH3_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] ch3_timer_rst_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                   // CH3_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> CH3_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          ch3_timer_rst_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                  // CH3_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> CH3_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          ch3_thresh_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                           // CH3_THRESH_s1_translator:uav_waitrequest -> CH3_THRESH_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] ch3_thresh_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                            // CH3_THRESH_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> CH3_THRESH_s1_translator:uav_burstcount
	wire   [31:0] ch3_thresh_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                             // CH3_THRESH_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> CH3_THRESH_s1_translator:uav_writedata
	wire   [21:0] ch3_thresh_s1_translator_avalon_universal_slave_0_agent_m0_address;                               // CH3_THRESH_s1_translator_avalon_universal_slave_0_agent:m0_address -> CH3_THRESH_s1_translator:uav_address
	wire          ch3_thresh_s1_translator_avalon_universal_slave_0_agent_m0_write;                                 // CH3_THRESH_s1_translator_avalon_universal_slave_0_agent:m0_write -> CH3_THRESH_s1_translator:uav_write
	wire          ch3_thresh_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                  // CH3_THRESH_s1_translator_avalon_universal_slave_0_agent:m0_lock -> CH3_THRESH_s1_translator:uav_lock
	wire          ch3_thresh_s1_translator_avalon_universal_slave_0_agent_m0_read;                                  // CH3_THRESH_s1_translator_avalon_universal_slave_0_agent:m0_read -> CH3_THRESH_s1_translator:uav_read
	wire   [31:0] ch3_thresh_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                              // CH3_THRESH_s1_translator:uav_readdata -> CH3_THRESH_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          ch3_thresh_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                         // CH3_THRESH_s1_translator:uav_readdatavalid -> CH3_THRESH_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          ch3_thresh_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                           // CH3_THRESH_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> CH3_THRESH_s1_translator:uav_debugaccess
	wire    [3:0] ch3_thresh_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                            // CH3_THRESH_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> CH3_THRESH_s1_translator:uav_byteenable
	wire          ch3_thresh_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                    // CH3_THRESH_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> CH3_THRESH_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          ch3_thresh_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                          // CH3_THRESH_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> CH3_THRESH_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          ch3_thresh_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                  // CH3_THRESH_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> CH3_THRESH_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] ch3_thresh_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                           // CH3_THRESH_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> CH3_THRESH_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          ch3_thresh_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                          // CH3_THRESH_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> CH3_THRESH_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          ch3_thresh_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                 // CH3_THRESH_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> CH3_THRESH_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          ch3_thresh_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                       // CH3_THRESH_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> CH3_THRESH_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          ch3_thresh_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;               // CH3_THRESH_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> CH3_THRESH_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] ch3_thresh_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                        // CH3_THRESH_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> CH3_THRESH_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          ch3_thresh_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                       // CH3_THRESH_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> CH3_THRESH_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          ch3_thresh_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                     // CH3_THRESH_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> CH3_THRESH_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] ch3_thresh_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                      // CH3_THRESH_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> CH3_THRESH_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          ch3_thresh_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                     // CH3_THRESH_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> CH3_THRESH_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          ch3_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                          // CH3_RD_PEAK_s1_translator:uav_waitrequest -> CH3_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] ch3_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                           // CH3_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> CH3_RD_PEAK_s1_translator:uav_burstcount
	wire   [31:0] ch3_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                            // CH3_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> CH3_RD_PEAK_s1_translator:uav_writedata
	wire   [21:0] ch3_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_address;                              // CH3_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:m0_address -> CH3_RD_PEAK_s1_translator:uav_address
	wire          ch3_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_write;                                // CH3_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:m0_write -> CH3_RD_PEAK_s1_translator:uav_write
	wire          ch3_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                 // CH3_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:m0_lock -> CH3_RD_PEAK_s1_translator:uav_lock
	wire          ch3_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_read;                                 // CH3_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:m0_read -> CH3_RD_PEAK_s1_translator:uav_read
	wire   [31:0] ch3_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                             // CH3_RD_PEAK_s1_translator:uav_readdata -> CH3_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          ch3_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                        // CH3_RD_PEAK_s1_translator:uav_readdatavalid -> CH3_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          ch3_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                          // CH3_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> CH3_RD_PEAK_s1_translator:uav_debugaccess
	wire    [3:0] ch3_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                           // CH3_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> CH3_RD_PEAK_s1_translator:uav_byteenable
	wire          ch3_rd_peak_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                   // CH3_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> CH3_RD_PEAK_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          ch3_rd_peak_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                         // CH3_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> CH3_RD_PEAK_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          ch3_rd_peak_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                 // CH3_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> CH3_RD_PEAK_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] ch3_rd_peak_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                          // CH3_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> CH3_RD_PEAK_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          ch3_rd_peak_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                         // CH3_RD_PEAK_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> CH3_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          ch3_rd_peak_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                // CH3_RD_PEAK_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> CH3_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          ch3_rd_peak_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                      // CH3_RD_PEAK_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> CH3_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          ch3_rd_peak_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;              // CH3_RD_PEAK_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> CH3_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] ch3_rd_peak_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                       // CH3_RD_PEAK_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> CH3_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          ch3_rd_peak_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                      // CH3_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> CH3_RD_PEAK_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          ch3_rd_peak_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                    // CH3_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> CH3_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] ch3_rd_peak_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                     // CH3_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> CH3_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          ch3_rd_peak_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                    // CH3_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> CH3_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          ch3_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                       // CH3_PEAK_FOUND_s1_translator:uav_waitrequest -> CH3_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] ch3_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                        // CH3_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> CH3_PEAK_FOUND_s1_translator:uav_burstcount
	wire   [31:0] ch3_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                         // CH3_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> CH3_PEAK_FOUND_s1_translator:uav_writedata
	wire   [21:0] ch3_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_address;                           // CH3_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:m0_address -> CH3_PEAK_FOUND_s1_translator:uav_address
	wire          ch3_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_write;                             // CH3_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:m0_write -> CH3_PEAK_FOUND_s1_translator:uav_write
	wire          ch3_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_lock;                              // CH3_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:m0_lock -> CH3_PEAK_FOUND_s1_translator:uav_lock
	wire          ch3_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_read;                              // CH3_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:m0_read -> CH3_PEAK_FOUND_s1_translator:uav_read
	wire   [31:0] ch3_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                          // CH3_PEAK_FOUND_s1_translator:uav_readdata -> CH3_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          ch3_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                     // CH3_PEAK_FOUND_s1_translator:uav_readdatavalid -> CH3_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          ch3_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                       // CH3_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> CH3_PEAK_FOUND_s1_translator:uav_debugaccess
	wire    [3:0] ch3_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                        // CH3_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> CH3_PEAK_FOUND_s1_translator:uav_byteenable
	wire          ch3_peak_found_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                // CH3_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> CH3_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          ch3_peak_found_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                      // CH3_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> CH3_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          ch3_peak_found_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;              // CH3_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> CH3_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] ch3_peak_found_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                       // CH3_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> CH3_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          ch3_peak_found_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                      // CH3_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> CH3_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          ch3_peak_found_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;             // CH3_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> CH3_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          ch3_peak_found_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                   // CH3_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> CH3_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          ch3_peak_found_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;           // CH3_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> CH3_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] ch3_peak_found_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                    // CH3_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> CH3_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          ch3_peak_found_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                   // CH3_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> CH3_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          ch3_peak_found_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                 // CH3_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> CH3_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] ch3_peak_found_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                  // CH3_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> CH3_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          ch3_peak_found_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                 // CH3_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> CH3_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          ch3_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                            // CH3_YN1_U_s1_translator:uav_waitrequest -> CH3_YN1_U_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] ch3_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                             // CH3_YN1_U_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> CH3_YN1_U_s1_translator:uav_burstcount
	wire   [31:0] ch3_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                              // CH3_YN1_U_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> CH3_YN1_U_s1_translator:uav_writedata
	wire   [21:0] ch3_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_address;                                // CH3_YN1_U_s1_translator_avalon_universal_slave_0_agent:m0_address -> CH3_YN1_U_s1_translator:uav_address
	wire          ch3_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_write;                                  // CH3_YN1_U_s1_translator_avalon_universal_slave_0_agent:m0_write -> CH3_YN1_U_s1_translator:uav_write
	wire          ch3_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                   // CH3_YN1_U_s1_translator_avalon_universal_slave_0_agent:m0_lock -> CH3_YN1_U_s1_translator:uav_lock
	wire          ch3_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_read;                                   // CH3_YN1_U_s1_translator_avalon_universal_slave_0_agent:m0_read -> CH3_YN1_U_s1_translator:uav_read
	wire   [31:0] ch3_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                               // CH3_YN1_U_s1_translator:uav_readdata -> CH3_YN1_U_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          ch3_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                          // CH3_YN1_U_s1_translator:uav_readdatavalid -> CH3_YN1_U_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          ch3_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                            // CH3_YN1_U_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> CH3_YN1_U_s1_translator:uav_debugaccess
	wire    [3:0] ch3_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                             // CH3_YN1_U_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> CH3_YN1_U_s1_translator:uav_byteenable
	wire          ch3_yn1_u_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                     // CH3_YN1_U_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> CH3_YN1_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          ch3_yn1_u_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                           // CH3_YN1_U_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> CH3_YN1_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          ch3_yn1_u_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                   // CH3_YN1_U_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> CH3_YN1_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] ch3_yn1_u_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                            // CH3_YN1_U_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> CH3_YN1_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          ch3_yn1_u_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                           // CH3_YN1_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> CH3_YN1_U_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          ch3_yn1_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                  // CH3_YN1_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> CH3_YN1_U_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          ch3_yn1_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                        // CH3_YN1_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> CH3_YN1_U_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          ch3_yn1_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                // CH3_YN1_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> CH3_YN1_U_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] ch3_yn1_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                         // CH3_YN1_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> CH3_YN1_U_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          ch3_yn1_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                        // CH3_YN1_U_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> CH3_YN1_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          ch3_yn1_u_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                      // CH3_YN1_U_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> CH3_YN1_U_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] ch3_yn1_u_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                       // CH3_YN1_U_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> CH3_YN1_U_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          ch3_yn1_u_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                      // CH3_YN1_U_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> CH3_YN1_U_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          ch3_time_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                             // CH3_TIME_s1_translator:uav_waitrequest -> CH3_TIME_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] ch3_time_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                              // CH3_TIME_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> CH3_TIME_s1_translator:uav_burstcount
	wire   [31:0] ch3_time_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                               // CH3_TIME_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> CH3_TIME_s1_translator:uav_writedata
	wire   [21:0] ch3_time_s1_translator_avalon_universal_slave_0_agent_m0_address;                                 // CH3_TIME_s1_translator_avalon_universal_slave_0_agent:m0_address -> CH3_TIME_s1_translator:uav_address
	wire          ch3_time_s1_translator_avalon_universal_slave_0_agent_m0_write;                                   // CH3_TIME_s1_translator_avalon_universal_slave_0_agent:m0_write -> CH3_TIME_s1_translator:uav_write
	wire          ch3_time_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                    // CH3_TIME_s1_translator_avalon_universal_slave_0_agent:m0_lock -> CH3_TIME_s1_translator:uav_lock
	wire          ch3_time_s1_translator_avalon_universal_slave_0_agent_m0_read;                                    // CH3_TIME_s1_translator_avalon_universal_slave_0_agent:m0_read -> CH3_TIME_s1_translator:uav_read
	wire   [31:0] ch3_time_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                // CH3_TIME_s1_translator:uav_readdata -> CH3_TIME_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          ch3_time_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                           // CH3_TIME_s1_translator:uav_readdatavalid -> CH3_TIME_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          ch3_time_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                             // CH3_TIME_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> CH3_TIME_s1_translator:uav_debugaccess
	wire    [3:0] ch3_time_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                              // CH3_TIME_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> CH3_TIME_s1_translator:uav_byteenable
	wire          ch3_time_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                      // CH3_TIME_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> CH3_TIME_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          ch3_time_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                            // CH3_TIME_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> CH3_TIME_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          ch3_time_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                    // CH3_TIME_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> CH3_TIME_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] ch3_time_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                             // CH3_TIME_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> CH3_TIME_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          ch3_time_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                            // CH3_TIME_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> CH3_TIME_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          ch3_time_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                   // CH3_TIME_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> CH3_TIME_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          ch3_time_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                         // CH3_TIME_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> CH3_TIME_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          ch3_time_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                 // CH3_TIME_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> CH3_TIME_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] ch3_time_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                          // CH3_TIME_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> CH3_TIME_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          ch3_time_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                         // CH3_TIME_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> CH3_TIME_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          ch3_time_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                       // CH3_TIME_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> CH3_TIME_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] ch3_time_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                        // CH3_TIME_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> CH3_TIME_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          ch3_time_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                       // CH3_TIME_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> CH3_TIME_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          ch3_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                            // CH3_YN3_L_s1_translator:uav_waitrequest -> CH3_YN3_L_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] ch3_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                             // CH3_YN3_L_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> CH3_YN3_L_s1_translator:uav_burstcount
	wire   [31:0] ch3_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                              // CH3_YN3_L_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> CH3_YN3_L_s1_translator:uav_writedata
	wire   [21:0] ch3_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_address;                                // CH3_YN3_L_s1_translator_avalon_universal_slave_0_agent:m0_address -> CH3_YN3_L_s1_translator:uav_address
	wire          ch3_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_write;                                  // CH3_YN3_L_s1_translator_avalon_universal_slave_0_agent:m0_write -> CH3_YN3_L_s1_translator:uav_write
	wire          ch3_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                   // CH3_YN3_L_s1_translator_avalon_universal_slave_0_agent:m0_lock -> CH3_YN3_L_s1_translator:uav_lock
	wire          ch3_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_read;                                   // CH3_YN3_L_s1_translator_avalon_universal_slave_0_agent:m0_read -> CH3_YN3_L_s1_translator:uav_read
	wire   [31:0] ch3_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                               // CH3_YN3_L_s1_translator:uav_readdata -> CH3_YN3_L_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          ch3_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                          // CH3_YN3_L_s1_translator:uav_readdatavalid -> CH3_YN3_L_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          ch3_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                            // CH3_YN3_L_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> CH3_YN3_L_s1_translator:uav_debugaccess
	wire    [3:0] ch3_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                             // CH3_YN3_L_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> CH3_YN3_L_s1_translator:uav_byteenable
	wire          ch3_yn3_l_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                     // CH3_YN3_L_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> CH3_YN3_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          ch3_yn3_l_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                           // CH3_YN3_L_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> CH3_YN3_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          ch3_yn3_l_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                   // CH3_YN3_L_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> CH3_YN3_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] ch3_yn3_l_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                            // CH3_YN3_L_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> CH3_YN3_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          ch3_yn3_l_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                           // CH3_YN3_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> CH3_YN3_L_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          ch3_yn3_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                  // CH3_YN3_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> CH3_YN3_L_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          ch3_yn3_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                        // CH3_YN3_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> CH3_YN3_L_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          ch3_yn3_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                // CH3_YN3_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> CH3_YN3_L_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] ch3_yn3_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                         // CH3_YN3_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> CH3_YN3_L_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          ch3_yn3_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                        // CH3_YN3_L_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> CH3_YN3_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          ch3_yn3_l_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                      // CH3_YN3_L_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> CH3_YN3_L_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] ch3_yn3_l_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                       // CH3_YN3_L_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> CH3_YN3_L_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          ch3_yn3_l_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                      // CH3_YN3_L_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> CH3_YN3_L_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          ch3_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                           // CH3_YN3_ML_s1_translator:uav_waitrequest -> CH3_YN3_ML_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] ch3_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                            // CH3_YN3_ML_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> CH3_YN3_ML_s1_translator:uav_burstcount
	wire   [31:0] ch3_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                             // CH3_YN3_ML_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> CH3_YN3_ML_s1_translator:uav_writedata
	wire   [21:0] ch3_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_address;                               // CH3_YN3_ML_s1_translator_avalon_universal_slave_0_agent:m0_address -> CH3_YN3_ML_s1_translator:uav_address
	wire          ch3_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_write;                                 // CH3_YN3_ML_s1_translator_avalon_universal_slave_0_agent:m0_write -> CH3_YN3_ML_s1_translator:uav_write
	wire          ch3_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                  // CH3_YN3_ML_s1_translator_avalon_universal_slave_0_agent:m0_lock -> CH3_YN3_ML_s1_translator:uav_lock
	wire          ch3_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_read;                                  // CH3_YN3_ML_s1_translator_avalon_universal_slave_0_agent:m0_read -> CH3_YN3_ML_s1_translator:uav_read
	wire   [31:0] ch3_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                              // CH3_YN3_ML_s1_translator:uav_readdata -> CH3_YN3_ML_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          ch3_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                         // CH3_YN3_ML_s1_translator:uav_readdatavalid -> CH3_YN3_ML_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          ch3_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                           // CH3_YN3_ML_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> CH3_YN3_ML_s1_translator:uav_debugaccess
	wire    [3:0] ch3_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                            // CH3_YN3_ML_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> CH3_YN3_ML_s1_translator:uav_byteenable
	wire          ch3_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                    // CH3_YN3_ML_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> CH3_YN3_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          ch3_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                          // CH3_YN3_ML_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> CH3_YN3_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          ch3_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                  // CH3_YN3_ML_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> CH3_YN3_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] ch3_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                           // CH3_YN3_ML_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> CH3_YN3_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          ch3_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                          // CH3_YN3_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> CH3_YN3_ML_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          ch3_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                 // CH3_YN3_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> CH3_YN3_ML_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          ch3_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                       // CH3_YN3_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> CH3_YN3_ML_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          ch3_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;               // CH3_YN3_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> CH3_YN3_ML_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] ch3_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                        // CH3_YN3_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> CH3_YN3_ML_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          ch3_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                       // CH3_YN3_ML_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> CH3_YN3_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          ch3_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                     // CH3_YN3_ML_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> CH3_YN3_ML_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] ch3_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                      // CH3_YN3_ML_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> CH3_YN3_ML_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          ch3_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                     // CH3_YN3_ML_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> CH3_YN3_ML_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          ch3_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                           // CH3_YN3_MU_s1_translator:uav_waitrequest -> CH3_YN3_MU_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] ch3_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                            // CH3_YN3_MU_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> CH3_YN3_MU_s1_translator:uav_burstcount
	wire   [31:0] ch3_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                             // CH3_YN3_MU_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> CH3_YN3_MU_s1_translator:uav_writedata
	wire   [21:0] ch3_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_address;                               // CH3_YN3_MU_s1_translator_avalon_universal_slave_0_agent:m0_address -> CH3_YN3_MU_s1_translator:uav_address
	wire          ch3_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_write;                                 // CH3_YN3_MU_s1_translator_avalon_universal_slave_0_agent:m0_write -> CH3_YN3_MU_s1_translator:uav_write
	wire          ch3_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                  // CH3_YN3_MU_s1_translator_avalon_universal_slave_0_agent:m0_lock -> CH3_YN3_MU_s1_translator:uav_lock
	wire          ch3_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_read;                                  // CH3_YN3_MU_s1_translator_avalon_universal_slave_0_agent:m0_read -> CH3_YN3_MU_s1_translator:uav_read
	wire   [31:0] ch3_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                              // CH3_YN3_MU_s1_translator:uav_readdata -> CH3_YN3_MU_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          ch3_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                         // CH3_YN3_MU_s1_translator:uav_readdatavalid -> CH3_YN3_MU_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          ch3_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                           // CH3_YN3_MU_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> CH3_YN3_MU_s1_translator:uav_debugaccess
	wire    [3:0] ch3_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                            // CH3_YN3_MU_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> CH3_YN3_MU_s1_translator:uav_byteenable
	wire          ch3_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                    // CH3_YN3_MU_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> CH3_YN3_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          ch3_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                          // CH3_YN3_MU_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> CH3_YN3_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          ch3_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                  // CH3_YN3_MU_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> CH3_YN3_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] ch3_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                           // CH3_YN3_MU_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> CH3_YN3_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          ch3_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                          // CH3_YN3_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> CH3_YN3_MU_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          ch3_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                 // CH3_YN3_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> CH3_YN3_MU_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          ch3_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                       // CH3_YN3_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> CH3_YN3_MU_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          ch3_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;               // CH3_YN3_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> CH3_YN3_MU_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] ch3_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                        // CH3_YN3_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> CH3_YN3_MU_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          ch3_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                       // CH3_YN3_MU_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> CH3_YN3_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          ch3_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                     // CH3_YN3_MU_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> CH3_YN3_MU_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] ch3_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                      // CH3_YN3_MU_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> CH3_YN3_MU_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          ch3_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                     // CH3_YN3_MU_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> CH3_YN3_MU_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          ch3_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                            // CH3_YN3_U_s1_translator:uav_waitrequest -> CH3_YN3_U_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] ch3_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                             // CH3_YN3_U_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> CH3_YN3_U_s1_translator:uav_burstcount
	wire   [31:0] ch3_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                              // CH3_YN3_U_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> CH3_YN3_U_s1_translator:uav_writedata
	wire   [21:0] ch3_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_address;                                // CH3_YN3_U_s1_translator_avalon_universal_slave_0_agent:m0_address -> CH3_YN3_U_s1_translator:uav_address
	wire          ch3_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_write;                                  // CH3_YN3_U_s1_translator_avalon_universal_slave_0_agent:m0_write -> CH3_YN3_U_s1_translator:uav_write
	wire          ch3_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                   // CH3_YN3_U_s1_translator_avalon_universal_slave_0_agent:m0_lock -> CH3_YN3_U_s1_translator:uav_lock
	wire          ch3_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_read;                                   // CH3_YN3_U_s1_translator_avalon_universal_slave_0_agent:m0_read -> CH3_YN3_U_s1_translator:uav_read
	wire   [31:0] ch3_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                               // CH3_YN3_U_s1_translator:uav_readdata -> CH3_YN3_U_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          ch3_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                          // CH3_YN3_U_s1_translator:uav_readdatavalid -> CH3_YN3_U_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          ch3_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                            // CH3_YN3_U_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> CH3_YN3_U_s1_translator:uav_debugaccess
	wire    [3:0] ch3_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                             // CH3_YN3_U_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> CH3_YN3_U_s1_translator:uav_byteenable
	wire          ch3_yn3_u_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                     // CH3_YN3_U_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> CH3_YN3_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          ch3_yn3_u_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                           // CH3_YN3_U_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> CH3_YN3_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          ch3_yn3_u_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                   // CH3_YN3_U_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> CH3_YN3_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] ch3_yn3_u_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                            // CH3_YN3_U_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> CH3_YN3_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          ch3_yn3_u_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                           // CH3_YN3_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> CH3_YN3_U_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          ch3_yn3_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                  // CH3_YN3_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> CH3_YN3_U_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          ch3_yn3_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                        // CH3_YN3_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> CH3_YN3_U_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          ch3_yn3_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                // CH3_YN3_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> CH3_YN3_U_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] ch3_yn3_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                         // CH3_YN3_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> CH3_YN3_U_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          ch3_yn3_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                        // CH3_YN3_U_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> CH3_YN3_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          ch3_yn3_u_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                      // CH3_YN3_U_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> CH3_YN3_U_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] ch3_yn3_u_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                       // CH3_YN3_U_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> CH3_YN3_U_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          ch3_yn3_u_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                      // CH3_YN3_U_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> CH3_YN3_U_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          ch3_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                            // CH3_YN2_L_s1_translator:uav_waitrequest -> CH3_YN2_L_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] ch3_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                             // CH3_YN2_L_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> CH3_YN2_L_s1_translator:uav_burstcount
	wire   [31:0] ch3_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                              // CH3_YN2_L_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> CH3_YN2_L_s1_translator:uav_writedata
	wire   [21:0] ch3_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_address;                                // CH3_YN2_L_s1_translator_avalon_universal_slave_0_agent:m0_address -> CH3_YN2_L_s1_translator:uav_address
	wire          ch3_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_write;                                  // CH3_YN2_L_s1_translator_avalon_universal_slave_0_agent:m0_write -> CH3_YN2_L_s1_translator:uav_write
	wire          ch3_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                   // CH3_YN2_L_s1_translator_avalon_universal_slave_0_agent:m0_lock -> CH3_YN2_L_s1_translator:uav_lock
	wire          ch3_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_read;                                   // CH3_YN2_L_s1_translator_avalon_universal_slave_0_agent:m0_read -> CH3_YN2_L_s1_translator:uav_read
	wire   [31:0] ch3_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                               // CH3_YN2_L_s1_translator:uav_readdata -> CH3_YN2_L_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          ch3_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                          // CH3_YN2_L_s1_translator:uav_readdatavalid -> CH3_YN2_L_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          ch3_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                            // CH3_YN2_L_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> CH3_YN2_L_s1_translator:uav_debugaccess
	wire    [3:0] ch3_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                             // CH3_YN2_L_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> CH3_YN2_L_s1_translator:uav_byteenable
	wire          ch3_yn2_l_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                     // CH3_YN2_L_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> CH3_YN2_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          ch3_yn2_l_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                           // CH3_YN2_L_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> CH3_YN2_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          ch3_yn2_l_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                   // CH3_YN2_L_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> CH3_YN2_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] ch3_yn2_l_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                            // CH3_YN2_L_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> CH3_YN2_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          ch3_yn2_l_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                           // CH3_YN2_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> CH3_YN2_L_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          ch3_yn2_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                  // CH3_YN2_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> CH3_YN2_L_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          ch3_yn2_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                        // CH3_YN2_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> CH3_YN2_L_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          ch3_yn2_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                // CH3_YN2_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> CH3_YN2_L_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] ch3_yn2_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                         // CH3_YN2_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> CH3_YN2_L_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          ch3_yn2_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                        // CH3_YN2_L_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> CH3_YN2_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          ch3_yn2_l_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                      // CH3_YN2_L_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> CH3_YN2_L_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] ch3_yn2_l_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                       // CH3_YN2_L_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> CH3_YN2_L_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          ch3_yn2_l_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                      // CH3_YN2_L_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> CH3_YN2_L_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          ch3_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                           // CH3_YN2_ML_s1_translator:uav_waitrequest -> CH3_YN2_ML_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] ch3_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                            // CH3_YN2_ML_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> CH3_YN2_ML_s1_translator:uav_burstcount
	wire   [31:0] ch3_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                             // CH3_YN2_ML_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> CH3_YN2_ML_s1_translator:uav_writedata
	wire   [21:0] ch3_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_address;                               // CH3_YN2_ML_s1_translator_avalon_universal_slave_0_agent:m0_address -> CH3_YN2_ML_s1_translator:uav_address
	wire          ch3_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_write;                                 // CH3_YN2_ML_s1_translator_avalon_universal_slave_0_agent:m0_write -> CH3_YN2_ML_s1_translator:uav_write
	wire          ch3_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                  // CH3_YN2_ML_s1_translator_avalon_universal_slave_0_agent:m0_lock -> CH3_YN2_ML_s1_translator:uav_lock
	wire          ch3_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_read;                                  // CH3_YN2_ML_s1_translator_avalon_universal_slave_0_agent:m0_read -> CH3_YN2_ML_s1_translator:uav_read
	wire   [31:0] ch3_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                              // CH3_YN2_ML_s1_translator:uav_readdata -> CH3_YN2_ML_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          ch3_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                         // CH3_YN2_ML_s1_translator:uav_readdatavalid -> CH3_YN2_ML_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          ch3_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                           // CH3_YN2_ML_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> CH3_YN2_ML_s1_translator:uav_debugaccess
	wire    [3:0] ch3_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                            // CH3_YN2_ML_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> CH3_YN2_ML_s1_translator:uav_byteenable
	wire          ch3_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                    // CH3_YN2_ML_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> CH3_YN2_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          ch3_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                          // CH3_YN2_ML_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> CH3_YN2_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          ch3_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                  // CH3_YN2_ML_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> CH3_YN2_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] ch3_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                           // CH3_YN2_ML_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> CH3_YN2_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          ch3_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                          // CH3_YN2_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> CH3_YN2_ML_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          ch3_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                 // CH3_YN2_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> CH3_YN2_ML_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          ch3_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                       // CH3_YN2_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> CH3_YN2_ML_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          ch3_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;               // CH3_YN2_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> CH3_YN2_ML_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] ch3_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                        // CH3_YN2_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> CH3_YN2_ML_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          ch3_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                       // CH3_YN2_ML_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> CH3_YN2_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          ch3_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                     // CH3_YN2_ML_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> CH3_YN2_ML_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] ch3_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                      // CH3_YN2_ML_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> CH3_YN2_ML_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          ch3_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                     // CH3_YN2_ML_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> CH3_YN2_ML_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          ch3_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                           // CH3_YN2_MU_s1_translator:uav_waitrequest -> CH3_YN2_MU_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] ch3_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                            // CH3_YN2_MU_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> CH3_YN2_MU_s1_translator:uav_burstcount
	wire   [31:0] ch3_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                             // CH3_YN2_MU_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> CH3_YN2_MU_s1_translator:uav_writedata
	wire   [21:0] ch3_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_address;                               // CH3_YN2_MU_s1_translator_avalon_universal_slave_0_agent:m0_address -> CH3_YN2_MU_s1_translator:uav_address
	wire          ch3_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_write;                                 // CH3_YN2_MU_s1_translator_avalon_universal_slave_0_agent:m0_write -> CH3_YN2_MU_s1_translator:uav_write
	wire          ch3_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                  // CH3_YN2_MU_s1_translator_avalon_universal_slave_0_agent:m0_lock -> CH3_YN2_MU_s1_translator:uav_lock
	wire          ch3_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_read;                                  // CH3_YN2_MU_s1_translator_avalon_universal_slave_0_agent:m0_read -> CH3_YN2_MU_s1_translator:uav_read
	wire   [31:0] ch3_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                              // CH3_YN2_MU_s1_translator:uav_readdata -> CH3_YN2_MU_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          ch3_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                         // CH3_YN2_MU_s1_translator:uav_readdatavalid -> CH3_YN2_MU_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          ch3_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                           // CH3_YN2_MU_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> CH3_YN2_MU_s1_translator:uav_debugaccess
	wire    [3:0] ch3_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                            // CH3_YN2_MU_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> CH3_YN2_MU_s1_translator:uav_byteenable
	wire          ch3_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                    // CH3_YN2_MU_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> CH3_YN2_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          ch3_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                          // CH3_YN2_MU_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> CH3_YN2_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          ch3_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                  // CH3_YN2_MU_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> CH3_YN2_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] ch3_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                           // CH3_YN2_MU_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> CH3_YN2_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          ch3_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                          // CH3_YN2_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> CH3_YN2_MU_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          ch3_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                 // CH3_YN2_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> CH3_YN2_MU_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          ch3_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                       // CH3_YN2_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> CH3_YN2_MU_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          ch3_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;               // CH3_YN2_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> CH3_YN2_MU_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] ch3_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                        // CH3_YN2_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> CH3_YN2_MU_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          ch3_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                       // CH3_YN2_MU_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> CH3_YN2_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          ch3_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                     // CH3_YN2_MU_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> CH3_YN2_MU_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] ch3_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                      // CH3_YN2_MU_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> CH3_YN2_MU_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          ch3_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                     // CH3_YN2_MU_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> CH3_YN2_MU_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          ch3_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                            // CH3_YN2_U_s1_translator:uav_waitrequest -> CH3_YN2_U_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] ch3_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                             // CH3_YN2_U_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> CH3_YN2_U_s1_translator:uav_burstcount
	wire   [31:0] ch3_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                              // CH3_YN2_U_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> CH3_YN2_U_s1_translator:uav_writedata
	wire   [21:0] ch3_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_address;                                // CH3_YN2_U_s1_translator_avalon_universal_slave_0_agent:m0_address -> CH3_YN2_U_s1_translator:uav_address
	wire          ch3_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_write;                                  // CH3_YN2_U_s1_translator_avalon_universal_slave_0_agent:m0_write -> CH3_YN2_U_s1_translator:uav_write
	wire          ch3_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                   // CH3_YN2_U_s1_translator_avalon_universal_slave_0_agent:m0_lock -> CH3_YN2_U_s1_translator:uav_lock
	wire          ch3_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_read;                                   // CH3_YN2_U_s1_translator_avalon_universal_slave_0_agent:m0_read -> CH3_YN2_U_s1_translator:uav_read
	wire   [31:0] ch3_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                               // CH3_YN2_U_s1_translator:uav_readdata -> CH3_YN2_U_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          ch3_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                          // CH3_YN2_U_s1_translator:uav_readdatavalid -> CH3_YN2_U_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          ch3_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                            // CH3_YN2_U_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> CH3_YN2_U_s1_translator:uav_debugaccess
	wire    [3:0] ch3_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                             // CH3_YN2_U_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> CH3_YN2_U_s1_translator:uav_byteenable
	wire          ch3_yn2_u_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                     // CH3_YN2_U_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> CH3_YN2_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          ch3_yn2_u_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                           // CH3_YN2_U_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> CH3_YN2_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          ch3_yn2_u_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                   // CH3_YN2_U_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> CH3_YN2_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] ch3_yn2_u_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                            // CH3_YN2_U_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> CH3_YN2_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          ch3_yn2_u_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                           // CH3_YN2_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> CH3_YN2_U_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          ch3_yn2_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                  // CH3_YN2_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> CH3_YN2_U_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          ch3_yn2_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                        // CH3_YN2_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> CH3_YN2_U_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          ch3_yn2_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                // CH3_YN2_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> CH3_YN2_U_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] ch3_yn2_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                         // CH3_YN2_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> CH3_YN2_U_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          ch3_yn2_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                        // CH3_YN2_U_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> CH3_YN2_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          ch3_yn2_u_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                      // CH3_YN2_U_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> CH3_YN2_U_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] ch3_yn2_u_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                       // CH3_YN2_U_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> CH3_YN2_U_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          ch3_yn2_u_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                      // CH3_YN2_U_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> CH3_YN2_U_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          ch3_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                            // CH3_YN1_L_s1_translator:uav_waitrequest -> CH3_YN1_L_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] ch3_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                             // CH3_YN1_L_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> CH3_YN1_L_s1_translator:uav_burstcount
	wire   [31:0] ch3_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                              // CH3_YN1_L_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> CH3_YN1_L_s1_translator:uav_writedata
	wire   [21:0] ch3_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_address;                                // CH3_YN1_L_s1_translator_avalon_universal_slave_0_agent:m0_address -> CH3_YN1_L_s1_translator:uav_address
	wire          ch3_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_write;                                  // CH3_YN1_L_s1_translator_avalon_universal_slave_0_agent:m0_write -> CH3_YN1_L_s1_translator:uav_write
	wire          ch3_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                   // CH3_YN1_L_s1_translator_avalon_universal_slave_0_agent:m0_lock -> CH3_YN1_L_s1_translator:uav_lock
	wire          ch3_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_read;                                   // CH3_YN1_L_s1_translator_avalon_universal_slave_0_agent:m0_read -> CH3_YN1_L_s1_translator:uav_read
	wire   [31:0] ch3_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                               // CH3_YN1_L_s1_translator:uav_readdata -> CH3_YN1_L_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          ch3_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                          // CH3_YN1_L_s1_translator:uav_readdatavalid -> CH3_YN1_L_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          ch3_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                            // CH3_YN1_L_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> CH3_YN1_L_s1_translator:uav_debugaccess
	wire    [3:0] ch3_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                             // CH3_YN1_L_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> CH3_YN1_L_s1_translator:uav_byteenable
	wire          ch3_yn1_l_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                     // CH3_YN1_L_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> CH3_YN1_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          ch3_yn1_l_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                           // CH3_YN1_L_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> CH3_YN1_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          ch3_yn1_l_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                   // CH3_YN1_L_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> CH3_YN1_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] ch3_yn1_l_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                            // CH3_YN1_L_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> CH3_YN1_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          ch3_yn1_l_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                           // CH3_YN1_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> CH3_YN1_L_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          ch3_yn1_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                  // CH3_YN1_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> CH3_YN1_L_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          ch3_yn1_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                        // CH3_YN1_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> CH3_YN1_L_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          ch3_yn1_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                // CH3_YN1_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> CH3_YN1_L_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] ch3_yn1_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                         // CH3_YN1_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> CH3_YN1_L_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          ch3_yn1_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                        // CH3_YN1_L_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> CH3_YN1_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          ch3_yn1_l_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                      // CH3_YN1_L_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> CH3_YN1_L_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] ch3_yn1_l_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                       // CH3_YN1_L_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> CH3_YN1_L_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          ch3_yn1_l_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                      // CH3_YN1_L_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> CH3_YN1_L_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          ch3_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                           // CH3_YN1_MU_s1_translator:uav_waitrequest -> CH3_YN1_MU_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] ch3_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                            // CH3_YN1_MU_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> CH3_YN1_MU_s1_translator:uav_burstcount
	wire   [31:0] ch3_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                             // CH3_YN1_MU_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> CH3_YN1_MU_s1_translator:uav_writedata
	wire   [21:0] ch3_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_address;                               // CH3_YN1_MU_s1_translator_avalon_universal_slave_0_agent:m0_address -> CH3_YN1_MU_s1_translator:uav_address
	wire          ch3_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_write;                                 // CH3_YN1_MU_s1_translator_avalon_universal_slave_0_agent:m0_write -> CH3_YN1_MU_s1_translator:uav_write
	wire          ch3_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                  // CH3_YN1_MU_s1_translator_avalon_universal_slave_0_agent:m0_lock -> CH3_YN1_MU_s1_translator:uav_lock
	wire          ch3_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_read;                                  // CH3_YN1_MU_s1_translator_avalon_universal_slave_0_agent:m0_read -> CH3_YN1_MU_s1_translator:uav_read
	wire   [31:0] ch3_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                              // CH3_YN1_MU_s1_translator:uav_readdata -> CH3_YN1_MU_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          ch3_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                         // CH3_YN1_MU_s1_translator:uav_readdatavalid -> CH3_YN1_MU_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          ch3_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                           // CH3_YN1_MU_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> CH3_YN1_MU_s1_translator:uav_debugaccess
	wire    [3:0] ch3_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                            // CH3_YN1_MU_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> CH3_YN1_MU_s1_translator:uav_byteenable
	wire          ch3_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                    // CH3_YN1_MU_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> CH3_YN1_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          ch3_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                          // CH3_YN1_MU_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> CH3_YN1_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          ch3_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                  // CH3_YN1_MU_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> CH3_YN1_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] ch3_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                           // CH3_YN1_MU_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> CH3_YN1_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          ch3_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                          // CH3_YN1_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> CH3_YN1_MU_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          ch3_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                 // CH3_YN1_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> CH3_YN1_MU_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          ch3_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                       // CH3_YN1_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> CH3_YN1_MU_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          ch3_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;               // CH3_YN1_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> CH3_YN1_MU_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] ch3_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                        // CH3_YN1_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> CH3_YN1_MU_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          ch3_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                       // CH3_YN1_MU_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> CH3_YN1_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          ch3_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                     // CH3_YN1_MU_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> CH3_YN1_MU_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] ch3_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                      // CH3_YN1_MU_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> CH3_YN1_MU_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          ch3_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                     // CH3_YN1_MU_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> CH3_YN1_MU_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          ch3_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                           // CH3_YN1_ML_s1_translator:uav_waitrequest -> CH3_YN1_ML_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] ch3_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                            // CH3_YN1_ML_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> CH3_YN1_ML_s1_translator:uav_burstcount
	wire   [31:0] ch3_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                             // CH3_YN1_ML_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> CH3_YN1_ML_s1_translator:uav_writedata
	wire   [21:0] ch3_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_address;                               // CH3_YN1_ML_s1_translator_avalon_universal_slave_0_agent:m0_address -> CH3_YN1_ML_s1_translator:uav_address
	wire          ch3_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_write;                                 // CH3_YN1_ML_s1_translator_avalon_universal_slave_0_agent:m0_write -> CH3_YN1_ML_s1_translator:uav_write
	wire          ch3_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                  // CH3_YN1_ML_s1_translator_avalon_universal_slave_0_agent:m0_lock -> CH3_YN1_ML_s1_translator:uav_lock
	wire          ch3_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_read;                                  // CH3_YN1_ML_s1_translator_avalon_universal_slave_0_agent:m0_read -> CH3_YN1_ML_s1_translator:uav_read
	wire   [31:0] ch3_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                              // CH3_YN1_ML_s1_translator:uav_readdata -> CH3_YN1_ML_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          ch3_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                         // CH3_YN1_ML_s1_translator:uav_readdatavalid -> CH3_YN1_ML_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          ch3_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                           // CH3_YN1_ML_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> CH3_YN1_ML_s1_translator:uav_debugaccess
	wire    [3:0] ch3_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                            // CH3_YN1_ML_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> CH3_YN1_ML_s1_translator:uav_byteenable
	wire          ch3_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                    // CH3_YN1_ML_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> CH3_YN1_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          ch3_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                          // CH3_YN1_ML_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> CH3_YN1_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          ch3_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                  // CH3_YN1_ML_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> CH3_YN1_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] ch3_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                           // CH3_YN1_ML_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> CH3_YN1_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          ch3_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                          // CH3_YN1_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> CH3_YN1_ML_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          ch3_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                 // CH3_YN1_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> CH3_YN1_ML_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          ch3_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                       // CH3_YN1_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> CH3_YN1_ML_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          ch3_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;               // CH3_YN1_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> CH3_YN1_ML_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] ch3_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                        // CH3_YN1_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> CH3_YN1_ML_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          ch3_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                       // CH3_YN1_ML_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> CH3_YN1_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          ch3_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                     // CH3_YN1_ML_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> CH3_YN1_ML_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] ch3_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                      // CH3_YN1_ML_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> CH3_YN1_ML_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          ch3_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                     // CH3_YN1_ML_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> CH3_YN1_ML_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          ch4_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                        // CH4_TIMER_RST_s1_translator:uav_waitrequest -> CH4_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] ch4_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                         // CH4_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> CH4_TIMER_RST_s1_translator:uav_burstcount
	wire   [31:0] ch4_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                          // CH4_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> CH4_TIMER_RST_s1_translator:uav_writedata
	wire   [21:0] ch4_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_address;                            // CH4_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:m0_address -> CH4_TIMER_RST_s1_translator:uav_address
	wire          ch4_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_write;                              // CH4_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:m0_write -> CH4_TIMER_RST_s1_translator:uav_write
	wire          ch4_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_lock;                               // CH4_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:m0_lock -> CH4_TIMER_RST_s1_translator:uav_lock
	wire          ch4_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_read;                               // CH4_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:m0_read -> CH4_TIMER_RST_s1_translator:uav_read
	wire   [31:0] ch4_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                           // CH4_TIMER_RST_s1_translator:uav_readdata -> CH4_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          ch4_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                      // CH4_TIMER_RST_s1_translator:uav_readdatavalid -> CH4_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          ch4_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                        // CH4_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> CH4_TIMER_RST_s1_translator:uav_debugaccess
	wire    [3:0] ch4_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                         // CH4_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> CH4_TIMER_RST_s1_translator:uav_byteenable
	wire          ch4_timer_rst_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                 // CH4_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> CH4_TIMER_RST_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          ch4_timer_rst_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                       // CH4_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> CH4_TIMER_RST_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          ch4_timer_rst_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;               // CH4_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> CH4_TIMER_RST_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] ch4_timer_rst_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                        // CH4_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> CH4_TIMER_RST_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          ch4_timer_rst_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                       // CH4_TIMER_RST_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> CH4_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          ch4_timer_rst_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;              // CH4_TIMER_RST_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> CH4_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          ch4_timer_rst_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                    // CH4_TIMER_RST_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> CH4_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          ch4_timer_rst_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;            // CH4_TIMER_RST_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> CH4_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] ch4_timer_rst_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                     // CH4_TIMER_RST_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> CH4_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          ch4_timer_rst_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                    // CH4_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> CH4_TIMER_RST_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          ch4_timer_rst_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                  // CH4_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> CH4_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] ch4_timer_rst_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                   // CH4_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> CH4_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          ch4_timer_rst_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                  // CH4_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> CH4_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          ch4_thresh_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                           // CH4_THRESH_s1_translator:uav_waitrequest -> CH4_THRESH_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] ch4_thresh_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                            // CH4_THRESH_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> CH4_THRESH_s1_translator:uav_burstcount
	wire   [31:0] ch4_thresh_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                             // CH4_THRESH_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> CH4_THRESH_s1_translator:uav_writedata
	wire   [21:0] ch4_thresh_s1_translator_avalon_universal_slave_0_agent_m0_address;                               // CH4_THRESH_s1_translator_avalon_universal_slave_0_agent:m0_address -> CH4_THRESH_s1_translator:uav_address
	wire          ch4_thresh_s1_translator_avalon_universal_slave_0_agent_m0_write;                                 // CH4_THRESH_s1_translator_avalon_universal_slave_0_agent:m0_write -> CH4_THRESH_s1_translator:uav_write
	wire          ch4_thresh_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                  // CH4_THRESH_s1_translator_avalon_universal_slave_0_agent:m0_lock -> CH4_THRESH_s1_translator:uav_lock
	wire          ch4_thresh_s1_translator_avalon_universal_slave_0_agent_m0_read;                                  // CH4_THRESH_s1_translator_avalon_universal_slave_0_agent:m0_read -> CH4_THRESH_s1_translator:uav_read
	wire   [31:0] ch4_thresh_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                              // CH4_THRESH_s1_translator:uav_readdata -> CH4_THRESH_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          ch4_thresh_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                         // CH4_THRESH_s1_translator:uav_readdatavalid -> CH4_THRESH_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          ch4_thresh_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                           // CH4_THRESH_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> CH4_THRESH_s1_translator:uav_debugaccess
	wire    [3:0] ch4_thresh_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                            // CH4_THRESH_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> CH4_THRESH_s1_translator:uav_byteenable
	wire          ch4_thresh_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                    // CH4_THRESH_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> CH4_THRESH_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          ch4_thresh_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                          // CH4_THRESH_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> CH4_THRESH_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          ch4_thresh_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                  // CH4_THRESH_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> CH4_THRESH_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] ch4_thresh_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                           // CH4_THRESH_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> CH4_THRESH_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          ch4_thresh_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                          // CH4_THRESH_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> CH4_THRESH_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          ch4_thresh_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                 // CH4_THRESH_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> CH4_THRESH_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          ch4_thresh_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                       // CH4_THRESH_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> CH4_THRESH_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          ch4_thresh_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;               // CH4_THRESH_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> CH4_THRESH_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] ch4_thresh_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                        // CH4_THRESH_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> CH4_THRESH_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          ch4_thresh_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                       // CH4_THRESH_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> CH4_THRESH_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          ch4_thresh_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                     // CH4_THRESH_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> CH4_THRESH_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] ch4_thresh_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                      // CH4_THRESH_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> CH4_THRESH_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          ch4_thresh_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                     // CH4_THRESH_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> CH4_THRESH_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          ch4_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                          // CH4_RD_PEAK_s1_translator:uav_waitrequest -> CH4_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] ch4_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                           // CH4_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> CH4_RD_PEAK_s1_translator:uav_burstcount
	wire   [31:0] ch4_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                            // CH4_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> CH4_RD_PEAK_s1_translator:uav_writedata
	wire   [21:0] ch4_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_address;                              // CH4_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:m0_address -> CH4_RD_PEAK_s1_translator:uav_address
	wire          ch4_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_write;                                // CH4_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:m0_write -> CH4_RD_PEAK_s1_translator:uav_write
	wire          ch4_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                 // CH4_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:m0_lock -> CH4_RD_PEAK_s1_translator:uav_lock
	wire          ch4_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_read;                                 // CH4_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:m0_read -> CH4_RD_PEAK_s1_translator:uav_read
	wire   [31:0] ch4_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                             // CH4_RD_PEAK_s1_translator:uav_readdata -> CH4_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          ch4_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                        // CH4_RD_PEAK_s1_translator:uav_readdatavalid -> CH4_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          ch4_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                          // CH4_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> CH4_RD_PEAK_s1_translator:uav_debugaccess
	wire    [3:0] ch4_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                           // CH4_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> CH4_RD_PEAK_s1_translator:uav_byteenable
	wire          ch4_rd_peak_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                   // CH4_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> CH4_RD_PEAK_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          ch4_rd_peak_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                         // CH4_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> CH4_RD_PEAK_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          ch4_rd_peak_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                 // CH4_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> CH4_RD_PEAK_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] ch4_rd_peak_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                          // CH4_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> CH4_RD_PEAK_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          ch4_rd_peak_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                         // CH4_RD_PEAK_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> CH4_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          ch4_rd_peak_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                // CH4_RD_PEAK_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> CH4_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          ch4_rd_peak_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                      // CH4_RD_PEAK_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> CH4_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          ch4_rd_peak_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;              // CH4_RD_PEAK_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> CH4_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] ch4_rd_peak_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                       // CH4_RD_PEAK_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> CH4_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          ch4_rd_peak_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                      // CH4_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> CH4_RD_PEAK_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          ch4_rd_peak_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                    // CH4_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> CH4_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] ch4_rd_peak_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                     // CH4_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> CH4_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          ch4_rd_peak_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                    // CH4_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> CH4_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          ch4_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                       // CH4_PEAK_FOUND_s1_translator:uav_waitrequest -> CH4_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] ch4_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                        // CH4_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> CH4_PEAK_FOUND_s1_translator:uav_burstcount
	wire   [31:0] ch4_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                         // CH4_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> CH4_PEAK_FOUND_s1_translator:uav_writedata
	wire   [21:0] ch4_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_address;                           // CH4_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:m0_address -> CH4_PEAK_FOUND_s1_translator:uav_address
	wire          ch4_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_write;                             // CH4_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:m0_write -> CH4_PEAK_FOUND_s1_translator:uav_write
	wire          ch4_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_lock;                              // CH4_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:m0_lock -> CH4_PEAK_FOUND_s1_translator:uav_lock
	wire          ch4_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_read;                              // CH4_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:m0_read -> CH4_PEAK_FOUND_s1_translator:uav_read
	wire   [31:0] ch4_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                          // CH4_PEAK_FOUND_s1_translator:uav_readdata -> CH4_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          ch4_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                     // CH4_PEAK_FOUND_s1_translator:uav_readdatavalid -> CH4_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          ch4_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                       // CH4_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> CH4_PEAK_FOUND_s1_translator:uav_debugaccess
	wire    [3:0] ch4_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                        // CH4_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> CH4_PEAK_FOUND_s1_translator:uav_byteenable
	wire          ch4_peak_found_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                // CH4_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> CH4_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          ch4_peak_found_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                      // CH4_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> CH4_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          ch4_peak_found_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;              // CH4_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> CH4_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] ch4_peak_found_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                       // CH4_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> CH4_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          ch4_peak_found_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                      // CH4_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> CH4_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          ch4_peak_found_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;             // CH4_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> CH4_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          ch4_peak_found_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                   // CH4_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> CH4_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          ch4_peak_found_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;           // CH4_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> CH4_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] ch4_peak_found_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                    // CH4_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> CH4_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          ch4_peak_found_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                   // CH4_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> CH4_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          ch4_peak_found_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                 // CH4_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> CH4_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] ch4_peak_found_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                  // CH4_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> CH4_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          ch4_peak_found_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                 // CH4_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> CH4_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          ch4_time_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                             // CH4_TIME_s1_translator:uav_waitrequest -> CH4_TIME_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] ch4_time_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                              // CH4_TIME_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> CH4_TIME_s1_translator:uav_burstcount
	wire   [31:0] ch4_time_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                               // CH4_TIME_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> CH4_TIME_s1_translator:uav_writedata
	wire   [21:0] ch4_time_s1_translator_avalon_universal_slave_0_agent_m0_address;                                 // CH4_TIME_s1_translator_avalon_universal_slave_0_agent:m0_address -> CH4_TIME_s1_translator:uav_address
	wire          ch4_time_s1_translator_avalon_universal_slave_0_agent_m0_write;                                   // CH4_TIME_s1_translator_avalon_universal_slave_0_agent:m0_write -> CH4_TIME_s1_translator:uav_write
	wire          ch4_time_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                    // CH4_TIME_s1_translator_avalon_universal_slave_0_agent:m0_lock -> CH4_TIME_s1_translator:uav_lock
	wire          ch4_time_s1_translator_avalon_universal_slave_0_agent_m0_read;                                    // CH4_TIME_s1_translator_avalon_universal_slave_0_agent:m0_read -> CH4_TIME_s1_translator:uav_read
	wire   [31:0] ch4_time_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                // CH4_TIME_s1_translator:uav_readdata -> CH4_TIME_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          ch4_time_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                           // CH4_TIME_s1_translator:uav_readdatavalid -> CH4_TIME_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          ch4_time_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                             // CH4_TIME_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> CH4_TIME_s1_translator:uav_debugaccess
	wire    [3:0] ch4_time_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                              // CH4_TIME_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> CH4_TIME_s1_translator:uav_byteenable
	wire          ch4_time_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                      // CH4_TIME_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> CH4_TIME_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          ch4_time_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                            // CH4_TIME_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> CH4_TIME_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          ch4_time_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                    // CH4_TIME_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> CH4_TIME_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] ch4_time_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                             // CH4_TIME_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> CH4_TIME_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          ch4_time_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                            // CH4_TIME_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> CH4_TIME_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          ch4_time_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                   // CH4_TIME_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> CH4_TIME_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          ch4_time_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                         // CH4_TIME_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> CH4_TIME_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          ch4_time_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                 // CH4_TIME_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> CH4_TIME_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] ch4_time_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                          // CH4_TIME_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> CH4_TIME_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          ch4_time_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                         // CH4_TIME_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> CH4_TIME_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          ch4_time_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                       // CH4_TIME_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> CH4_TIME_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] ch4_time_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                        // CH4_TIME_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> CH4_TIME_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          ch4_time_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                       // CH4_TIME_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> CH4_TIME_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          ch4_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                            // CH4_YN1_U_s1_translator:uav_waitrequest -> CH4_YN1_U_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] ch4_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                             // CH4_YN1_U_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> CH4_YN1_U_s1_translator:uav_burstcount
	wire   [31:0] ch4_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                              // CH4_YN1_U_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> CH4_YN1_U_s1_translator:uav_writedata
	wire   [21:0] ch4_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_address;                                // CH4_YN1_U_s1_translator_avalon_universal_slave_0_agent:m0_address -> CH4_YN1_U_s1_translator:uav_address
	wire          ch4_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_write;                                  // CH4_YN1_U_s1_translator_avalon_universal_slave_0_agent:m0_write -> CH4_YN1_U_s1_translator:uav_write
	wire          ch4_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                   // CH4_YN1_U_s1_translator_avalon_universal_slave_0_agent:m0_lock -> CH4_YN1_U_s1_translator:uav_lock
	wire          ch4_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_read;                                   // CH4_YN1_U_s1_translator_avalon_universal_slave_0_agent:m0_read -> CH4_YN1_U_s1_translator:uav_read
	wire   [31:0] ch4_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                               // CH4_YN1_U_s1_translator:uav_readdata -> CH4_YN1_U_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          ch4_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                          // CH4_YN1_U_s1_translator:uav_readdatavalid -> CH4_YN1_U_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          ch4_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                            // CH4_YN1_U_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> CH4_YN1_U_s1_translator:uav_debugaccess
	wire    [3:0] ch4_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                             // CH4_YN1_U_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> CH4_YN1_U_s1_translator:uav_byteenable
	wire          ch4_yn1_u_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                     // CH4_YN1_U_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> CH4_YN1_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          ch4_yn1_u_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                           // CH4_YN1_U_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> CH4_YN1_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          ch4_yn1_u_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                   // CH4_YN1_U_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> CH4_YN1_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] ch4_yn1_u_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                            // CH4_YN1_U_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> CH4_YN1_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          ch4_yn1_u_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                           // CH4_YN1_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> CH4_YN1_U_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          ch4_yn1_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                  // CH4_YN1_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> CH4_YN1_U_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          ch4_yn1_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                        // CH4_YN1_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> CH4_YN1_U_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          ch4_yn1_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                // CH4_YN1_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> CH4_YN1_U_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] ch4_yn1_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                         // CH4_YN1_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> CH4_YN1_U_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          ch4_yn1_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                        // CH4_YN1_U_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> CH4_YN1_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          ch4_yn1_u_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                      // CH4_YN1_U_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> CH4_YN1_U_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] ch4_yn1_u_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                       // CH4_YN1_U_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> CH4_YN1_U_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          ch4_yn1_u_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                      // CH4_YN1_U_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> CH4_YN1_U_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          ch4_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                           // CH4_YN1_MU_s1_translator:uav_waitrequest -> CH4_YN1_MU_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] ch4_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                            // CH4_YN1_MU_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> CH4_YN1_MU_s1_translator:uav_burstcount
	wire   [31:0] ch4_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                             // CH4_YN1_MU_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> CH4_YN1_MU_s1_translator:uav_writedata
	wire   [21:0] ch4_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_address;                               // CH4_YN1_MU_s1_translator_avalon_universal_slave_0_agent:m0_address -> CH4_YN1_MU_s1_translator:uav_address
	wire          ch4_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_write;                                 // CH4_YN1_MU_s1_translator_avalon_universal_slave_0_agent:m0_write -> CH4_YN1_MU_s1_translator:uav_write
	wire          ch4_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                  // CH4_YN1_MU_s1_translator_avalon_universal_slave_0_agent:m0_lock -> CH4_YN1_MU_s1_translator:uav_lock
	wire          ch4_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_read;                                  // CH4_YN1_MU_s1_translator_avalon_universal_slave_0_agent:m0_read -> CH4_YN1_MU_s1_translator:uav_read
	wire   [31:0] ch4_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                              // CH4_YN1_MU_s1_translator:uav_readdata -> CH4_YN1_MU_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          ch4_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                         // CH4_YN1_MU_s1_translator:uav_readdatavalid -> CH4_YN1_MU_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          ch4_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                           // CH4_YN1_MU_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> CH4_YN1_MU_s1_translator:uav_debugaccess
	wire    [3:0] ch4_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                            // CH4_YN1_MU_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> CH4_YN1_MU_s1_translator:uav_byteenable
	wire          ch4_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                    // CH4_YN1_MU_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> CH4_YN1_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          ch4_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                          // CH4_YN1_MU_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> CH4_YN1_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          ch4_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                  // CH4_YN1_MU_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> CH4_YN1_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] ch4_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                           // CH4_YN1_MU_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> CH4_YN1_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          ch4_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                          // CH4_YN1_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> CH4_YN1_MU_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          ch4_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                 // CH4_YN1_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> CH4_YN1_MU_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          ch4_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                       // CH4_YN1_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> CH4_YN1_MU_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          ch4_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;               // CH4_YN1_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> CH4_YN1_MU_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] ch4_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                        // CH4_YN1_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> CH4_YN1_MU_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          ch4_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                       // CH4_YN1_MU_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> CH4_YN1_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          ch4_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                     // CH4_YN1_MU_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> CH4_YN1_MU_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] ch4_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                      // CH4_YN1_MU_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> CH4_YN1_MU_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          ch4_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                     // CH4_YN1_MU_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> CH4_YN1_MU_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          ch4_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                           // CH4_YN1_ML_s1_translator:uav_waitrequest -> CH4_YN1_ML_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] ch4_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                            // CH4_YN1_ML_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> CH4_YN1_ML_s1_translator:uav_burstcount
	wire   [31:0] ch4_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                             // CH4_YN1_ML_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> CH4_YN1_ML_s1_translator:uav_writedata
	wire   [21:0] ch4_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_address;                               // CH4_YN1_ML_s1_translator_avalon_universal_slave_0_agent:m0_address -> CH4_YN1_ML_s1_translator:uav_address
	wire          ch4_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_write;                                 // CH4_YN1_ML_s1_translator_avalon_universal_slave_0_agent:m0_write -> CH4_YN1_ML_s1_translator:uav_write
	wire          ch4_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                  // CH4_YN1_ML_s1_translator_avalon_universal_slave_0_agent:m0_lock -> CH4_YN1_ML_s1_translator:uav_lock
	wire          ch4_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_read;                                  // CH4_YN1_ML_s1_translator_avalon_universal_slave_0_agent:m0_read -> CH4_YN1_ML_s1_translator:uav_read
	wire   [31:0] ch4_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                              // CH4_YN1_ML_s1_translator:uav_readdata -> CH4_YN1_ML_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          ch4_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                         // CH4_YN1_ML_s1_translator:uav_readdatavalid -> CH4_YN1_ML_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          ch4_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                           // CH4_YN1_ML_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> CH4_YN1_ML_s1_translator:uav_debugaccess
	wire    [3:0] ch4_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                            // CH4_YN1_ML_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> CH4_YN1_ML_s1_translator:uav_byteenable
	wire          ch4_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                    // CH4_YN1_ML_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> CH4_YN1_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          ch4_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                          // CH4_YN1_ML_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> CH4_YN1_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          ch4_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                  // CH4_YN1_ML_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> CH4_YN1_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] ch4_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                           // CH4_YN1_ML_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> CH4_YN1_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          ch4_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                          // CH4_YN1_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> CH4_YN1_ML_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          ch4_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                 // CH4_YN1_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> CH4_YN1_ML_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          ch4_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                       // CH4_YN1_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> CH4_YN1_ML_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          ch4_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;               // CH4_YN1_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> CH4_YN1_ML_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] ch4_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                        // CH4_YN1_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> CH4_YN1_ML_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          ch4_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                       // CH4_YN1_ML_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> CH4_YN1_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          ch4_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                     // CH4_YN1_ML_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> CH4_YN1_ML_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] ch4_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                      // CH4_YN1_ML_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> CH4_YN1_ML_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          ch4_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                     // CH4_YN1_ML_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> CH4_YN1_ML_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          ch4_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                            // CH4_YN1_L_s1_translator:uav_waitrequest -> CH4_YN1_L_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] ch4_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                             // CH4_YN1_L_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> CH4_YN1_L_s1_translator:uav_burstcount
	wire   [31:0] ch4_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                              // CH4_YN1_L_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> CH4_YN1_L_s1_translator:uav_writedata
	wire   [21:0] ch4_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_address;                                // CH4_YN1_L_s1_translator_avalon_universal_slave_0_agent:m0_address -> CH4_YN1_L_s1_translator:uav_address
	wire          ch4_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_write;                                  // CH4_YN1_L_s1_translator_avalon_universal_slave_0_agent:m0_write -> CH4_YN1_L_s1_translator:uav_write
	wire          ch4_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                   // CH4_YN1_L_s1_translator_avalon_universal_slave_0_agent:m0_lock -> CH4_YN1_L_s1_translator:uav_lock
	wire          ch4_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_read;                                   // CH4_YN1_L_s1_translator_avalon_universal_slave_0_agent:m0_read -> CH4_YN1_L_s1_translator:uav_read
	wire   [31:0] ch4_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                               // CH4_YN1_L_s1_translator:uav_readdata -> CH4_YN1_L_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          ch4_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                          // CH4_YN1_L_s1_translator:uav_readdatavalid -> CH4_YN1_L_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          ch4_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                            // CH4_YN1_L_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> CH4_YN1_L_s1_translator:uav_debugaccess
	wire    [3:0] ch4_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                             // CH4_YN1_L_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> CH4_YN1_L_s1_translator:uav_byteenable
	wire          ch4_yn1_l_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                     // CH4_YN1_L_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> CH4_YN1_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          ch4_yn1_l_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                           // CH4_YN1_L_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> CH4_YN1_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          ch4_yn1_l_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                   // CH4_YN1_L_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> CH4_YN1_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] ch4_yn1_l_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                            // CH4_YN1_L_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> CH4_YN1_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          ch4_yn1_l_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                           // CH4_YN1_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> CH4_YN1_L_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          ch4_yn1_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                  // CH4_YN1_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> CH4_YN1_L_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          ch4_yn1_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                        // CH4_YN1_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> CH4_YN1_L_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          ch4_yn1_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                // CH4_YN1_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> CH4_YN1_L_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] ch4_yn1_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                         // CH4_YN1_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> CH4_YN1_L_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          ch4_yn1_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                        // CH4_YN1_L_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> CH4_YN1_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          ch4_yn1_l_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                      // CH4_YN1_L_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> CH4_YN1_L_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] ch4_yn1_l_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                       // CH4_YN1_L_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> CH4_YN1_L_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          ch4_yn1_l_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                      // CH4_YN1_L_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> CH4_YN1_L_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          ch4_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                            // CH4_YN2_U_s1_translator:uav_waitrequest -> CH4_YN2_U_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] ch4_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                             // CH4_YN2_U_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> CH4_YN2_U_s1_translator:uav_burstcount
	wire   [31:0] ch4_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                              // CH4_YN2_U_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> CH4_YN2_U_s1_translator:uav_writedata
	wire   [21:0] ch4_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_address;                                // CH4_YN2_U_s1_translator_avalon_universal_slave_0_agent:m0_address -> CH4_YN2_U_s1_translator:uav_address
	wire          ch4_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_write;                                  // CH4_YN2_U_s1_translator_avalon_universal_slave_0_agent:m0_write -> CH4_YN2_U_s1_translator:uav_write
	wire          ch4_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                   // CH4_YN2_U_s1_translator_avalon_universal_slave_0_agent:m0_lock -> CH4_YN2_U_s1_translator:uav_lock
	wire          ch4_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_read;                                   // CH4_YN2_U_s1_translator_avalon_universal_slave_0_agent:m0_read -> CH4_YN2_U_s1_translator:uav_read
	wire   [31:0] ch4_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                               // CH4_YN2_U_s1_translator:uav_readdata -> CH4_YN2_U_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          ch4_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                          // CH4_YN2_U_s1_translator:uav_readdatavalid -> CH4_YN2_U_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          ch4_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                            // CH4_YN2_U_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> CH4_YN2_U_s1_translator:uav_debugaccess
	wire    [3:0] ch4_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                             // CH4_YN2_U_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> CH4_YN2_U_s1_translator:uav_byteenable
	wire          ch4_yn2_u_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                     // CH4_YN2_U_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> CH4_YN2_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          ch4_yn2_u_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                           // CH4_YN2_U_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> CH4_YN2_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          ch4_yn2_u_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                   // CH4_YN2_U_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> CH4_YN2_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] ch4_yn2_u_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                            // CH4_YN2_U_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> CH4_YN2_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          ch4_yn2_u_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                           // CH4_YN2_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> CH4_YN2_U_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          ch4_yn2_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                  // CH4_YN2_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> CH4_YN2_U_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          ch4_yn2_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                        // CH4_YN2_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> CH4_YN2_U_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          ch4_yn2_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                // CH4_YN2_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> CH4_YN2_U_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] ch4_yn2_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                         // CH4_YN2_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> CH4_YN2_U_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          ch4_yn2_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                        // CH4_YN2_U_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> CH4_YN2_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          ch4_yn2_u_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                      // CH4_YN2_U_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> CH4_YN2_U_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] ch4_yn2_u_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                       // CH4_YN2_U_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> CH4_YN2_U_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          ch4_yn2_u_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                      // CH4_YN2_U_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> CH4_YN2_U_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          ch4_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                           // CH4_YN2_MU_s1_translator:uav_waitrequest -> CH4_YN2_MU_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] ch4_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                            // CH4_YN2_MU_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> CH4_YN2_MU_s1_translator:uav_burstcount
	wire   [31:0] ch4_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                             // CH4_YN2_MU_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> CH4_YN2_MU_s1_translator:uav_writedata
	wire   [21:0] ch4_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_address;                               // CH4_YN2_MU_s1_translator_avalon_universal_slave_0_agent:m0_address -> CH4_YN2_MU_s1_translator:uav_address
	wire          ch4_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_write;                                 // CH4_YN2_MU_s1_translator_avalon_universal_slave_0_agent:m0_write -> CH4_YN2_MU_s1_translator:uav_write
	wire          ch4_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                  // CH4_YN2_MU_s1_translator_avalon_universal_slave_0_agent:m0_lock -> CH4_YN2_MU_s1_translator:uav_lock
	wire          ch4_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_read;                                  // CH4_YN2_MU_s1_translator_avalon_universal_slave_0_agent:m0_read -> CH4_YN2_MU_s1_translator:uav_read
	wire   [31:0] ch4_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                              // CH4_YN2_MU_s1_translator:uav_readdata -> CH4_YN2_MU_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          ch4_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                         // CH4_YN2_MU_s1_translator:uav_readdatavalid -> CH4_YN2_MU_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          ch4_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                           // CH4_YN2_MU_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> CH4_YN2_MU_s1_translator:uav_debugaccess
	wire    [3:0] ch4_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                            // CH4_YN2_MU_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> CH4_YN2_MU_s1_translator:uav_byteenable
	wire          ch4_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                    // CH4_YN2_MU_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> CH4_YN2_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          ch4_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                          // CH4_YN2_MU_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> CH4_YN2_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          ch4_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                  // CH4_YN2_MU_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> CH4_YN2_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] ch4_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                           // CH4_YN2_MU_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> CH4_YN2_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          ch4_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                          // CH4_YN2_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> CH4_YN2_MU_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          ch4_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                 // CH4_YN2_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> CH4_YN2_MU_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          ch4_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                       // CH4_YN2_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> CH4_YN2_MU_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          ch4_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;               // CH4_YN2_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> CH4_YN2_MU_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] ch4_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                        // CH4_YN2_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> CH4_YN2_MU_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          ch4_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                       // CH4_YN2_MU_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> CH4_YN2_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          ch4_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                     // CH4_YN2_MU_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> CH4_YN2_MU_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] ch4_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                      // CH4_YN2_MU_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> CH4_YN2_MU_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          ch4_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                     // CH4_YN2_MU_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> CH4_YN2_MU_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          ch4_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                           // CH4_YN2_ML_s1_translator:uav_waitrequest -> CH4_YN2_ML_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] ch4_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                            // CH4_YN2_ML_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> CH4_YN2_ML_s1_translator:uav_burstcount
	wire   [31:0] ch4_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                             // CH4_YN2_ML_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> CH4_YN2_ML_s1_translator:uav_writedata
	wire   [21:0] ch4_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_address;                               // CH4_YN2_ML_s1_translator_avalon_universal_slave_0_agent:m0_address -> CH4_YN2_ML_s1_translator:uav_address
	wire          ch4_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_write;                                 // CH4_YN2_ML_s1_translator_avalon_universal_slave_0_agent:m0_write -> CH4_YN2_ML_s1_translator:uav_write
	wire          ch4_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                  // CH4_YN2_ML_s1_translator_avalon_universal_slave_0_agent:m0_lock -> CH4_YN2_ML_s1_translator:uav_lock
	wire          ch4_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_read;                                  // CH4_YN2_ML_s1_translator_avalon_universal_slave_0_agent:m0_read -> CH4_YN2_ML_s1_translator:uav_read
	wire   [31:0] ch4_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                              // CH4_YN2_ML_s1_translator:uav_readdata -> CH4_YN2_ML_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          ch4_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                         // CH4_YN2_ML_s1_translator:uav_readdatavalid -> CH4_YN2_ML_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          ch4_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                           // CH4_YN2_ML_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> CH4_YN2_ML_s1_translator:uav_debugaccess
	wire    [3:0] ch4_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                            // CH4_YN2_ML_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> CH4_YN2_ML_s1_translator:uav_byteenable
	wire          ch4_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                    // CH4_YN2_ML_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> CH4_YN2_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          ch4_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                          // CH4_YN2_ML_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> CH4_YN2_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          ch4_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                  // CH4_YN2_ML_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> CH4_YN2_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] ch4_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                           // CH4_YN2_ML_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> CH4_YN2_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          ch4_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                          // CH4_YN2_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> CH4_YN2_ML_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          ch4_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                 // CH4_YN2_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> CH4_YN2_ML_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          ch4_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                       // CH4_YN2_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> CH4_YN2_ML_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          ch4_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;               // CH4_YN2_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> CH4_YN2_ML_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] ch4_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                        // CH4_YN2_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> CH4_YN2_ML_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          ch4_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                       // CH4_YN2_ML_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> CH4_YN2_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          ch4_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                     // CH4_YN2_ML_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> CH4_YN2_ML_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] ch4_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                      // CH4_YN2_ML_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> CH4_YN2_ML_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          ch4_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                     // CH4_YN2_ML_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> CH4_YN2_ML_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          ch4_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                            // CH4_YN2_L_s1_translator:uav_waitrequest -> CH4_YN2_L_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] ch4_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                             // CH4_YN2_L_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> CH4_YN2_L_s1_translator:uav_burstcount
	wire   [31:0] ch4_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                              // CH4_YN2_L_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> CH4_YN2_L_s1_translator:uav_writedata
	wire   [21:0] ch4_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_address;                                // CH4_YN2_L_s1_translator_avalon_universal_slave_0_agent:m0_address -> CH4_YN2_L_s1_translator:uav_address
	wire          ch4_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_write;                                  // CH4_YN2_L_s1_translator_avalon_universal_slave_0_agent:m0_write -> CH4_YN2_L_s1_translator:uav_write
	wire          ch4_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                   // CH4_YN2_L_s1_translator_avalon_universal_slave_0_agent:m0_lock -> CH4_YN2_L_s1_translator:uav_lock
	wire          ch4_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_read;                                   // CH4_YN2_L_s1_translator_avalon_universal_slave_0_agent:m0_read -> CH4_YN2_L_s1_translator:uav_read
	wire   [31:0] ch4_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                               // CH4_YN2_L_s1_translator:uav_readdata -> CH4_YN2_L_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          ch4_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                          // CH4_YN2_L_s1_translator:uav_readdatavalid -> CH4_YN2_L_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          ch4_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                            // CH4_YN2_L_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> CH4_YN2_L_s1_translator:uav_debugaccess
	wire    [3:0] ch4_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                             // CH4_YN2_L_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> CH4_YN2_L_s1_translator:uav_byteenable
	wire          ch4_yn2_l_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                     // CH4_YN2_L_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> CH4_YN2_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          ch4_yn2_l_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                           // CH4_YN2_L_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> CH4_YN2_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          ch4_yn2_l_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                   // CH4_YN2_L_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> CH4_YN2_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] ch4_yn2_l_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                            // CH4_YN2_L_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> CH4_YN2_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          ch4_yn2_l_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                           // CH4_YN2_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> CH4_YN2_L_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          ch4_yn2_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                  // CH4_YN2_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> CH4_YN2_L_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          ch4_yn2_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                        // CH4_YN2_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> CH4_YN2_L_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          ch4_yn2_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                // CH4_YN2_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> CH4_YN2_L_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] ch4_yn2_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                         // CH4_YN2_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> CH4_YN2_L_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          ch4_yn2_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                        // CH4_YN2_L_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> CH4_YN2_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          ch4_yn2_l_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                      // CH4_YN2_L_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> CH4_YN2_L_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] ch4_yn2_l_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                       // CH4_YN2_L_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> CH4_YN2_L_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          ch4_yn2_l_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                      // CH4_YN2_L_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> CH4_YN2_L_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          ch4_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                            // CH4_YN3_U_s1_translator:uav_waitrequest -> CH4_YN3_U_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] ch4_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                             // CH4_YN3_U_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> CH4_YN3_U_s1_translator:uav_burstcount
	wire   [31:0] ch4_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                              // CH4_YN3_U_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> CH4_YN3_U_s1_translator:uav_writedata
	wire   [21:0] ch4_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_address;                                // CH4_YN3_U_s1_translator_avalon_universal_slave_0_agent:m0_address -> CH4_YN3_U_s1_translator:uav_address
	wire          ch4_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_write;                                  // CH4_YN3_U_s1_translator_avalon_universal_slave_0_agent:m0_write -> CH4_YN3_U_s1_translator:uav_write
	wire          ch4_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                   // CH4_YN3_U_s1_translator_avalon_universal_slave_0_agent:m0_lock -> CH4_YN3_U_s1_translator:uav_lock
	wire          ch4_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_read;                                   // CH4_YN3_U_s1_translator_avalon_universal_slave_0_agent:m0_read -> CH4_YN3_U_s1_translator:uav_read
	wire   [31:0] ch4_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                               // CH4_YN3_U_s1_translator:uav_readdata -> CH4_YN3_U_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          ch4_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                          // CH4_YN3_U_s1_translator:uav_readdatavalid -> CH4_YN3_U_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          ch4_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                            // CH4_YN3_U_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> CH4_YN3_U_s1_translator:uav_debugaccess
	wire    [3:0] ch4_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                             // CH4_YN3_U_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> CH4_YN3_U_s1_translator:uav_byteenable
	wire          ch4_yn3_u_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                     // CH4_YN3_U_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> CH4_YN3_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          ch4_yn3_u_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                           // CH4_YN3_U_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> CH4_YN3_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          ch4_yn3_u_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                   // CH4_YN3_U_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> CH4_YN3_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] ch4_yn3_u_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                            // CH4_YN3_U_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> CH4_YN3_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          ch4_yn3_u_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                           // CH4_YN3_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> CH4_YN3_U_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          ch4_yn3_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                  // CH4_YN3_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> CH4_YN3_U_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          ch4_yn3_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                        // CH4_YN3_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> CH4_YN3_U_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          ch4_yn3_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                // CH4_YN3_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> CH4_YN3_U_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] ch4_yn3_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                         // CH4_YN3_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> CH4_YN3_U_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          ch4_yn3_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                        // CH4_YN3_U_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> CH4_YN3_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          ch4_yn3_u_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                      // CH4_YN3_U_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> CH4_YN3_U_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] ch4_yn3_u_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                       // CH4_YN3_U_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> CH4_YN3_U_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          ch4_yn3_u_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                      // CH4_YN3_U_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> CH4_YN3_U_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          ch4_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                           // CH4_YN3_MU_s1_translator:uav_waitrequest -> CH4_YN3_MU_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] ch4_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                            // CH4_YN3_MU_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> CH4_YN3_MU_s1_translator:uav_burstcount
	wire   [31:0] ch4_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                             // CH4_YN3_MU_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> CH4_YN3_MU_s1_translator:uav_writedata
	wire   [21:0] ch4_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_address;                               // CH4_YN3_MU_s1_translator_avalon_universal_slave_0_agent:m0_address -> CH4_YN3_MU_s1_translator:uav_address
	wire          ch4_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_write;                                 // CH4_YN3_MU_s1_translator_avalon_universal_slave_0_agent:m0_write -> CH4_YN3_MU_s1_translator:uav_write
	wire          ch4_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                  // CH4_YN3_MU_s1_translator_avalon_universal_slave_0_agent:m0_lock -> CH4_YN3_MU_s1_translator:uav_lock
	wire          ch4_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_read;                                  // CH4_YN3_MU_s1_translator_avalon_universal_slave_0_agent:m0_read -> CH4_YN3_MU_s1_translator:uav_read
	wire   [31:0] ch4_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                              // CH4_YN3_MU_s1_translator:uav_readdata -> CH4_YN3_MU_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          ch4_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                         // CH4_YN3_MU_s1_translator:uav_readdatavalid -> CH4_YN3_MU_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          ch4_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                           // CH4_YN3_MU_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> CH4_YN3_MU_s1_translator:uav_debugaccess
	wire    [3:0] ch4_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                            // CH4_YN3_MU_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> CH4_YN3_MU_s1_translator:uav_byteenable
	wire          ch4_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                    // CH4_YN3_MU_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> CH4_YN3_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          ch4_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                          // CH4_YN3_MU_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> CH4_YN3_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          ch4_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                  // CH4_YN3_MU_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> CH4_YN3_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] ch4_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                           // CH4_YN3_MU_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> CH4_YN3_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          ch4_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                          // CH4_YN3_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> CH4_YN3_MU_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          ch4_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                 // CH4_YN3_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> CH4_YN3_MU_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          ch4_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                       // CH4_YN3_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> CH4_YN3_MU_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          ch4_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;               // CH4_YN3_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> CH4_YN3_MU_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] ch4_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                        // CH4_YN3_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> CH4_YN3_MU_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          ch4_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                       // CH4_YN3_MU_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> CH4_YN3_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          ch4_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                     // CH4_YN3_MU_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> CH4_YN3_MU_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] ch4_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                      // CH4_YN3_MU_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> CH4_YN3_MU_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          ch4_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                     // CH4_YN3_MU_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> CH4_YN3_MU_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          ch4_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                           // CH4_YN3_ML_s1_translator:uav_waitrequest -> CH4_YN3_ML_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] ch4_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                            // CH4_YN3_ML_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> CH4_YN3_ML_s1_translator:uav_burstcount
	wire   [31:0] ch4_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                             // CH4_YN3_ML_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> CH4_YN3_ML_s1_translator:uav_writedata
	wire   [21:0] ch4_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_address;                               // CH4_YN3_ML_s1_translator_avalon_universal_slave_0_agent:m0_address -> CH4_YN3_ML_s1_translator:uav_address
	wire          ch4_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_write;                                 // CH4_YN3_ML_s1_translator_avalon_universal_slave_0_agent:m0_write -> CH4_YN3_ML_s1_translator:uav_write
	wire          ch4_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                  // CH4_YN3_ML_s1_translator_avalon_universal_slave_0_agent:m0_lock -> CH4_YN3_ML_s1_translator:uav_lock
	wire          ch4_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_read;                                  // CH4_YN3_ML_s1_translator_avalon_universal_slave_0_agent:m0_read -> CH4_YN3_ML_s1_translator:uav_read
	wire   [31:0] ch4_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                              // CH4_YN3_ML_s1_translator:uav_readdata -> CH4_YN3_ML_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          ch4_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                         // CH4_YN3_ML_s1_translator:uav_readdatavalid -> CH4_YN3_ML_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          ch4_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                           // CH4_YN3_ML_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> CH4_YN3_ML_s1_translator:uav_debugaccess
	wire    [3:0] ch4_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                            // CH4_YN3_ML_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> CH4_YN3_ML_s1_translator:uav_byteenable
	wire          ch4_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                    // CH4_YN3_ML_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> CH4_YN3_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          ch4_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                          // CH4_YN3_ML_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> CH4_YN3_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          ch4_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                  // CH4_YN3_ML_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> CH4_YN3_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] ch4_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                           // CH4_YN3_ML_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> CH4_YN3_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          ch4_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                          // CH4_YN3_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> CH4_YN3_ML_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          ch4_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                 // CH4_YN3_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> CH4_YN3_ML_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          ch4_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                       // CH4_YN3_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> CH4_YN3_ML_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          ch4_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;               // CH4_YN3_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> CH4_YN3_ML_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] ch4_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                        // CH4_YN3_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> CH4_YN3_ML_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          ch4_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                       // CH4_YN3_ML_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> CH4_YN3_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          ch4_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                     // CH4_YN3_ML_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> CH4_YN3_ML_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] ch4_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                      // CH4_YN3_ML_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> CH4_YN3_ML_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          ch4_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                     // CH4_YN3_ML_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> CH4_YN3_ML_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          ch4_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                            // CH4_YN3_L_s1_translator:uav_waitrequest -> CH4_YN3_L_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] ch4_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                             // CH4_YN3_L_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> CH4_YN3_L_s1_translator:uav_burstcount
	wire   [31:0] ch4_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                              // CH4_YN3_L_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> CH4_YN3_L_s1_translator:uav_writedata
	wire   [21:0] ch4_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_address;                                // CH4_YN3_L_s1_translator_avalon_universal_slave_0_agent:m0_address -> CH4_YN3_L_s1_translator:uav_address
	wire          ch4_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_write;                                  // CH4_YN3_L_s1_translator_avalon_universal_slave_0_agent:m0_write -> CH4_YN3_L_s1_translator:uav_write
	wire          ch4_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                   // CH4_YN3_L_s1_translator_avalon_universal_slave_0_agent:m0_lock -> CH4_YN3_L_s1_translator:uav_lock
	wire          ch4_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_read;                                   // CH4_YN3_L_s1_translator_avalon_universal_slave_0_agent:m0_read -> CH4_YN3_L_s1_translator:uav_read
	wire   [31:0] ch4_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                               // CH4_YN3_L_s1_translator:uav_readdata -> CH4_YN3_L_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          ch4_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                          // CH4_YN3_L_s1_translator:uav_readdatavalid -> CH4_YN3_L_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          ch4_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                            // CH4_YN3_L_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> CH4_YN3_L_s1_translator:uav_debugaccess
	wire    [3:0] ch4_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                             // CH4_YN3_L_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> CH4_YN3_L_s1_translator:uav_byteenable
	wire          ch4_yn3_l_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                     // CH4_YN3_L_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> CH4_YN3_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          ch4_yn3_l_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                           // CH4_YN3_L_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> CH4_YN3_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          ch4_yn3_l_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                   // CH4_YN3_L_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> CH4_YN3_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] ch4_yn3_l_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                            // CH4_YN3_L_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> CH4_YN3_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          ch4_yn3_l_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                           // CH4_YN3_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> CH4_YN3_L_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          ch4_yn3_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                  // CH4_YN3_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> CH4_YN3_L_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          ch4_yn3_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                        // CH4_YN3_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> CH4_YN3_L_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          ch4_yn3_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                // CH4_YN3_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> CH4_YN3_L_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] ch4_yn3_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                         // CH4_YN3_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> CH4_YN3_L_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          ch4_yn3_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                        // CH4_YN3_L_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> CH4_YN3_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          ch4_yn3_l_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                      // CH4_YN3_L_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> CH4_YN3_L_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] ch4_yn3_l_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                       // CH4_YN3_L_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> CH4_YN3_L_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          ch4_yn3_l_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                      // CH4_YN3_L_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> CH4_YN3_L_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          nios_cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket;            // NIOS_CPU_instruction_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router:sink_endofpacket
	wire          nios_cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_valid;                  // NIOS_CPU_instruction_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router:sink_valid
	wire          nios_cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket;          // NIOS_CPU_instruction_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router:sink_startofpacket
	wire  [102:0] nios_cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_data;                   // NIOS_CPU_instruction_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router:sink_data
	wire          nios_cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_ready;                  // addr_router:sink_ready -> NIOS_CPU_instruction_master_translator_avalon_universal_master_0_agent:cp_ready
	wire          nios_cpu_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                   // NIOS_CPU_data_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_001:sink_endofpacket
	wire          nios_cpu_data_master_translator_avalon_universal_master_0_agent_cp_valid;                         // NIOS_CPU_data_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_001:sink_valid
	wire          nios_cpu_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket;                 // NIOS_CPU_data_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_001:sink_startofpacket
	wire  [102:0] nios_cpu_data_master_translator_avalon_universal_master_0_agent_cp_data;                          // NIOS_CPU_data_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_001:sink_data
	wire          nios_cpu_data_master_translator_avalon_universal_master_0_agent_cp_ready;                         // addr_router_001:sink_ready -> NIOS_CPU_data_master_translator_avalon_universal_master_0_agent:cp_ready
	wire          nios_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket;              // NIOS_CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router:sink_endofpacket
	wire          nios_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid;                    // NIOS_CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_valid -> id_router:sink_valid
	wire          nios_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket;            // NIOS_CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router:sink_startofpacket
	wire  [102:0] nios_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data;                     // NIOS_CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_data -> id_router:sink_data
	wire          nios_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready;                    // id_router:sink_ready -> NIOS_CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_ready
	wire          ram_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                  // RAM_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_001:sink_endofpacket
	wire          ram_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                        // RAM_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_001:sink_valid
	wire          ram_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                // RAM_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_001:sink_startofpacket
	wire  [102:0] ram_s1_translator_avalon_universal_slave_0_agent_rp_data;                                         // RAM_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_001:sink_data
	wire          ram_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                        // id_router_001:sink_ready -> RAM_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          ssram_uas_translator_avalon_universal_slave_0_agent_rp_endofpacket;                               // SSRAM_uas_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_002:sink_endofpacket
	wire          ssram_uas_translator_avalon_universal_slave_0_agent_rp_valid;                                     // SSRAM_uas_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_002:sink_valid
	wire          ssram_uas_translator_avalon_universal_slave_0_agent_rp_startofpacket;                             // SSRAM_uas_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_002:sink_startofpacket
	wire  [102:0] ssram_uas_translator_avalon_universal_slave_0_agent_rp_data;                                      // SSRAM_uas_translator_avalon_universal_slave_0_agent:rp_data -> id_router_002:sink_data
	wire          ssram_uas_translator_avalon_universal_slave_0_agent_rp_ready;                                     // id_router_002:sink_ready -> SSRAM_uas_translator_avalon_universal_slave_0_agent:rp_ready
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;             // JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_003:sink_endofpacket
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid;                   // JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_003:sink_valid
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;           // JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_003:sink_startofpacket
	wire  [102:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data;                    // JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_003:sink_data
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready;                   // id_router_003:sink_ready -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          lcd_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                       // LCD_control_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_004:sink_endofpacket
	wire          lcd_control_slave_translator_avalon_universal_slave_0_agent_rp_valid;                             // LCD_control_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_004:sink_valid
	wire          lcd_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                     // LCD_control_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_004:sink_startofpacket
	wire  [102:0] lcd_control_slave_translator_avalon_universal_slave_0_agent_rp_data;                              // LCD_control_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_004:sink_data
	wire          lcd_control_slave_translator_avalon_universal_slave_0_agent_rp_ready;                             // id_router_004:sink_ready -> LCD_control_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          adc_on_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                               // ADC_ON_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_005:sink_endofpacket
	wire          adc_on_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                     // ADC_ON_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_005:sink_valid
	wire          adc_on_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                             // ADC_ON_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_005:sink_startofpacket
	wire  [102:0] adc_on_s1_translator_avalon_universal_slave_0_agent_rp_data;                                      // ADC_ON_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_005:sink_data
	wire          adc_on_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                     // id_router_005:sink_ready -> ADC_ON_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          fifo_adc_data_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                        // FIFO_ADC_DATA_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_006:sink_endofpacket
	wire          fifo_adc_data_s1_translator_avalon_universal_slave_0_agent_rp_valid;                              // FIFO_ADC_DATA_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_006:sink_valid
	wire          fifo_adc_data_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                      // FIFO_ADC_DATA_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_006:sink_startofpacket
	wire  [102:0] fifo_adc_data_s1_translator_avalon_universal_slave_0_agent_rp_data;                               // FIFO_ADC_DATA_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_006:sink_data
	wire          fifo_adc_data_s1_translator_avalon_universal_slave_0_agent_rp_ready;                              // id_router_006:sink_ready -> FIFO_ADC_DATA_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          fifo_adc_data_valid_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                  // FIFO_ADC_DATA_VALID_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_007:sink_endofpacket
	wire          fifo_adc_data_valid_s1_translator_avalon_universal_slave_0_agent_rp_valid;                        // FIFO_ADC_DATA_VALID_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_007:sink_valid
	wire          fifo_adc_data_valid_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                // FIFO_ADC_DATA_VALID_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_007:sink_startofpacket
	wire  [102:0] fifo_adc_data_valid_s1_translator_avalon_universal_slave_0_agent_rp_data;                         // FIFO_ADC_DATA_VALID_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_007:sink_data
	wire          fifo_adc_data_valid_s1_translator_avalon_universal_slave_0_agent_rp_ready;                        // id_router_007:sink_ready -> FIFO_ADC_DATA_VALID_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          fifo_rst_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                             // FIFO_RST_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_008:sink_endofpacket
	wire          fifo_rst_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                   // FIFO_RST_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_008:sink_valid
	wire          fifo_rst_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                           // FIFO_RST_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_008:sink_startofpacket
	wire  [102:0] fifo_rst_s1_translator_avalon_universal_slave_0_agent_rp_data;                                    // FIFO_RST_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_008:sink_data
	wire          fifo_rst_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                   // id_router_008:sink_ready -> FIFO_RST_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          subtractor_on_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                        // SUBTRACTOR_ON_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_009:sink_endofpacket
	wire          subtractor_on_s1_translator_avalon_universal_slave_0_agent_rp_valid;                              // SUBTRACTOR_ON_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_009:sink_valid
	wire          subtractor_on_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                      // SUBTRACTOR_ON_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_009:sink_startofpacket
	wire  [102:0] subtractor_on_s1_translator_avalon_universal_slave_0_agent_rp_data;                               // SUBTRACTOR_ON_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_009:sink_data
	wire          subtractor_on_s1_translator_avalon_universal_slave_0_agent_rp_ready;                              // id_router_009:sink_ready -> SUBTRACTOR_ON_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          ch0_timer_rst_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                        // CH0_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_010:sink_endofpacket
	wire          ch0_timer_rst_s1_translator_avalon_universal_slave_0_agent_rp_valid;                              // CH0_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_010:sink_valid
	wire          ch0_timer_rst_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                      // CH0_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_010:sink_startofpacket
	wire  [102:0] ch0_timer_rst_s1_translator_avalon_universal_slave_0_agent_rp_data;                               // CH0_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_010:sink_data
	wire          ch0_timer_rst_s1_translator_avalon_universal_slave_0_agent_rp_ready;                              // id_router_010:sink_ready -> CH0_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          detector_on_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                          // DETECTOR_ON_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_011:sink_endofpacket
	wire          detector_on_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                // DETECTOR_ON_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_011:sink_valid
	wire          detector_on_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                        // DETECTOR_ON_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_011:sink_startofpacket
	wire  [102:0] detector_on_s1_translator_avalon_universal_slave_0_agent_rp_data;                                 // DETECTOR_ON_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_011:sink_data
	wire          detector_on_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                // id_router_011:sink_ready -> DETECTOR_ON_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          menu_down_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                            // MENU_DOWN_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_012:sink_endofpacket
	wire          menu_down_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                  // MENU_DOWN_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_012:sink_valid
	wire          menu_down_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                          // MENU_DOWN_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_012:sink_startofpacket
	wire  [102:0] menu_down_s1_translator_avalon_universal_slave_0_agent_rp_data;                                   // MENU_DOWN_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_012:sink_data
	wire          menu_down_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                  // id_router_012:sink_ready -> MENU_DOWN_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          menu_up_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                              // MENU_UP_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_013:sink_endofpacket
	wire          menu_up_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                    // MENU_UP_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_013:sink_valid
	wire          menu_up_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                            // MENU_UP_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_013:sink_startofpacket
	wire  [102:0] menu_up_s1_translator_avalon_universal_slave_0_agent_rp_data;                                     // MENU_UP_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_013:sink_data
	wire          menu_up_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                    // id_router_013:sink_ready -> MENU_UP_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          menu_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                 // MENU_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_014:sink_endofpacket
	wire          menu_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                       // MENU_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_014:sink_valid
	wire          menu_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                               // MENU_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_014:sink_startofpacket
	wire  [102:0] menu_s1_translator_avalon_universal_slave_0_agent_rp_data;                                        // MENU_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_014:sink_data
	wire          menu_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                       // id_router_014:sink_ready -> MENU_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          ch0_thresh_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                           // CH0_THRESH_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_015:sink_endofpacket
	wire          ch0_thresh_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                 // CH0_THRESH_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_015:sink_valid
	wire          ch0_thresh_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                         // CH0_THRESH_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_015:sink_startofpacket
	wire  [102:0] ch0_thresh_s1_translator_avalon_universal_slave_0_agent_rp_data;                                  // CH0_THRESH_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_015:sink_data
	wire          ch0_thresh_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                 // id_router_015:sink_ready -> CH0_THRESH_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          ch0_rd_peak_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                          // CH0_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_016:sink_endofpacket
	wire          ch0_rd_peak_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                // CH0_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_016:sink_valid
	wire          ch0_rd_peak_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                        // CH0_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_016:sink_startofpacket
	wire  [102:0] ch0_rd_peak_s1_translator_avalon_universal_slave_0_agent_rp_data;                                 // CH0_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_016:sink_data
	wire          ch0_rd_peak_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                // id_router_016:sink_ready -> CH0_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          ch0_peak_found_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                       // CH0_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_017:sink_endofpacket
	wire          ch0_peak_found_s1_translator_avalon_universal_slave_0_agent_rp_valid;                             // CH0_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_017:sink_valid
	wire          ch0_peak_found_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                     // CH0_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_017:sink_startofpacket
	wire  [102:0] ch0_peak_found_s1_translator_avalon_universal_slave_0_agent_rp_data;                              // CH0_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_017:sink_data
	wire          ch0_peak_found_s1_translator_avalon_universal_slave_0_agent_rp_ready;                             // id_router_017:sink_ready -> CH0_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          ch0_yn1_l_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                            // CH0_YN1_L_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_018:sink_endofpacket
	wire          ch0_yn1_l_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                  // CH0_YN1_L_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_018:sink_valid
	wire          ch0_yn1_l_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                          // CH0_YN1_L_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_018:sink_startofpacket
	wire  [102:0] ch0_yn1_l_s1_translator_avalon_universal_slave_0_agent_rp_data;                                   // CH0_YN1_L_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_018:sink_data
	wire          ch0_yn1_l_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                  // id_router_018:sink_ready -> CH0_YN1_L_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          ch0_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                           // CH0_YN1_ML_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_019:sink_endofpacket
	wire          ch0_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                 // CH0_YN1_ML_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_019:sink_valid
	wire          ch0_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                         // CH0_YN1_ML_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_019:sink_startofpacket
	wire  [102:0] ch0_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rp_data;                                  // CH0_YN1_ML_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_019:sink_data
	wire          ch0_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                 // id_router_019:sink_ready -> CH0_YN1_ML_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          ch0_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                           // CH0_YN1_MU_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_020:sink_endofpacket
	wire          ch0_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                 // CH0_YN1_MU_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_020:sink_valid
	wire          ch0_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                         // CH0_YN1_MU_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_020:sink_startofpacket
	wire  [102:0] ch0_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rp_data;                                  // CH0_YN1_MU_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_020:sink_data
	wire          ch0_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                 // id_router_020:sink_ready -> CH0_YN1_MU_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          ch0_yn1_u_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                            // CH0_YN1_U_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_021:sink_endofpacket
	wire          ch0_yn1_u_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                  // CH0_YN1_U_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_021:sink_valid
	wire          ch0_yn1_u_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                          // CH0_YN1_U_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_021:sink_startofpacket
	wire  [102:0] ch0_yn1_u_s1_translator_avalon_universal_slave_0_agent_rp_data;                                   // CH0_YN1_U_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_021:sink_data
	wire          ch0_yn1_u_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                  // id_router_021:sink_ready -> CH0_YN1_U_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          ch0_time_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                             // CH0_TIME_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_022:sink_endofpacket
	wire          ch0_time_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                   // CH0_TIME_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_022:sink_valid
	wire          ch0_time_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                           // CH0_TIME_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_022:sink_startofpacket
	wire  [102:0] ch0_time_s1_translator_avalon_universal_slave_0_agent_rp_data;                                    // CH0_TIME_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_022:sink_data
	wire          ch0_time_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                   // id_router_022:sink_ready -> CH0_TIME_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          ch0_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                           // CH0_YN2_MU_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_023:sink_endofpacket
	wire          ch0_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                 // CH0_YN2_MU_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_023:sink_valid
	wire          ch0_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                         // CH0_YN2_MU_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_023:sink_startofpacket
	wire  [102:0] ch0_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rp_data;                                  // CH0_YN2_MU_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_023:sink_data
	wire          ch0_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                 // id_router_023:sink_ready -> CH0_YN2_MU_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          ch0_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                           // CH0_YN2_ML_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_024:sink_endofpacket
	wire          ch0_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                 // CH0_YN2_ML_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_024:sink_valid
	wire          ch0_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                         // CH0_YN2_ML_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_024:sink_startofpacket
	wire  [102:0] ch0_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rp_data;                                  // CH0_YN2_ML_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_024:sink_data
	wire          ch0_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                 // id_router_024:sink_ready -> CH0_YN2_ML_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          ch0_yn2_u_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                            // CH0_YN2_U_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_025:sink_endofpacket
	wire          ch0_yn2_u_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                  // CH0_YN2_U_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_025:sink_valid
	wire          ch0_yn2_u_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                          // CH0_YN2_U_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_025:sink_startofpacket
	wire  [102:0] ch0_yn2_u_s1_translator_avalon_universal_slave_0_agent_rp_data;                                   // CH0_YN2_U_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_025:sink_data
	wire          ch0_yn2_u_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                  // id_router_025:sink_ready -> CH0_YN2_U_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          ch0_yn2_l_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                            // CH0_YN2_L_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_026:sink_endofpacket
	wire          ch0_yn2_l_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                  // CH0_YN2_L_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_026:sink_valid
	wire          ch0_yn2_l_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                          // CH0_YN2_L_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_026:sink_startofpacket
	wire  [102:0] ch0_yn2_l_s1_translator_avalon_universal_slave_0_agent_rp_data;                                   // CH0_YN2_L_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_026:sink_data
	wire          ch0_yn2_l_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                  // id_router_026:sink_ready -> CH0_YN2_L_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          ch0_yn3_l_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                            // CH0_YN3_L_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_027:sink_endofpacket
	wire          ch0_yn3_l_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                  // CH0_YN3_L_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_027:sink_valid
	wire          ch0_yn3_l_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                          // CH0_YN3_L_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_027:sink_startofpacket
	wire  [102:0] ch0_yn3_l_s1_translator_avalon_universal_slave_0_agent_rp_data;                                   // CH0_YN3_L_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_027:sink_data
	wire          ch0_yn3_l_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                  // id_router_027:sink_ready -> CH0_YN3_L_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          ch0_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                           // CH0_YN3_ML_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_028:sink_endofpacket
	wire          ch0_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                 // CH0_YN3_ML_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_028:sink_valid
	wire          ch0_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                         // CH0_YN3_ML_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_028:sink_startofpacket
	wire  [102:0] ch0_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rp_data;                                  // CH0_YN3_ML_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_028:sink_data
	wire          ch0_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                 // id_router_028:sink_ready -> CH0_YN3_ML_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          ch0_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                           // CH0_YN3_MU_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_029:sink_endofpacket
	wire          ch0_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                 // CH0_YN3_MU_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_029:sink_valid
	wire          ch0_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                         // CH0_YN3_MU_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_029:sink_startofpacket
	wire  [102:0] ch0_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rp_data;                                  // CH0_YN3_MU_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_029:sink_data
	wire          ch0_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                 // id_router_029:sink_ready -> CH0_YN3_MU_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          ch0_yn3_u_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                            // CH0_YN3_U_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_030:sink_endofpacket
	wire          ch0_yn3_u_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                  // CH0_YN3_U_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_030:sink_valid
	wire          ch0_yn3_u_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                          // CH0_YN3_U_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_030:sink_startofpacket
	wire  [102:0] ch0_yn3_u_s1_translator_avalon_universal_slave_0_agent_rp_data;                                   // CH0_YN3_U_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_030:sink_data
	wire          ch0_yn3_u_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                  // id_router_030:sink_ready -> CH0_YN3_U_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          ch1_timer_rst_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                        // CH1_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_031:sink_endofpacket
	wire          ch1_timer_rst_s1_translator_avalon_universal_slave_0_agent_rp_valid;                              // CH1_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_031:sink_valid
	wire          ch1_timer_rst_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                      // CH1_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_031:sink_startofpacket
	wire  [102:0] ch1_timer_rst_s1_translator_avalon_universal_slave_0_agent_rp_data;                               // CH1_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_031:sink_data
	wire          ch1_timer_rst_s1_translator_avalon_universal_slave_0_agent_rp_ready;                              // id_router_031:sink_ready -> CH1_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          ch1_thresh_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                           // CH1_THRESH_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_032:sink_endofpacket
	wire          ch1_thresh_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                 // CH1_THRESH_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_032:sink_valid
	wire          ch1_thresh_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                         // CH1_THRESH_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_032:sink_startofpacket
	wire  [102:0] ch1_thresh_s1_translator_avalon_universal_slave_0_agent_rp_data;                                  // CH1_THRESH_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_032:sink_data
	wire          ch1_thresh_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                 // id_router_032:sink_ready -> CH1_THRESH_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          ch1_rd_peak_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                          // CH1_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_033:sink_endofpacket
	wire          ch1_rd_peak_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                // CH1_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_033:sink_valid
	wire          ch1_rd_peak_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                        // CH1_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_033:sink_startofpacket
	wire  [102:0] ch1_rd_peak_s1_translator_avalon_universal_slave_0_agent_rp_data;                                 // CH1_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_033:sink_data
	wire          ch1_rd_peak_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                // id_router_033:sink_ready -> CH1_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          ch1_peak_found_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                       // CH1_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_034:sink_endofpacket
	wire          ch1_peak_found_s1_translator_avalon_universal_slave_0_agent_rp_valid;                             // CH1_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_034:sink_valid
	wire          ch1_peak_found_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                     // CH1_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_034:sink_startofpacket
	wire  [102:0] ch1_peak_found_s1_translator_avalon_universal_slave_0_agent_rp_data;                              // CH1_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_034:sink_data
	wire          ch1_peak_found_s1_translator_avalon_universal_slave_0_agent_rp_ready;                             // id_router_034:sink_ready -> CH1_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          ch1_time_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                             // CH1_TIME_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_035:sink_endofpacket
	wire          ch1_time_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                   // CH1_TIME_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_035:sink_valid
	wire          ch1_time_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                           // CH1_TIME_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_035:sink_startofpacket
	wire  [102:0] ch1_time_s1_translator_avalon_universal_slave_0_agent_rp_data;                                    // CH1_TIME_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_035:sink_data
	wire          ch1_time_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                   // id_router_035:sink_ready -> CH1_TIME_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          ch1_yn1_u_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                            // CH1_YN1_U_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_036:sink_endofpacket
	wire          ch1_yn1_u_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                  // CH1_YN1_U_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_036:sink_valid
	wire          ch1_yn1_u_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                          // CH1_YN1_U_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_036:sink_startofpacket
	wire  [102:0] ch1_yn1_u_s1_translator_avalon_universal_slave_0_agent_rp_data;                                   // CH1_YN1_U_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_036:sink_data
	wire          ch1_yn1_u_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                  // id_router_036:sink_ready -> CH1_YN1_U_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          ch1_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                           // CH1_YN1_MU_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_037:sink_endofpacket
	wire          ch1_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                 // CH1_YN1_MU_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_037:sink_valid
	wire          ch1_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                         // CH1_YN1_MU_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_037:sink_startofpacket
	wire  [102:0] ch1_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rp_data;                                  // CH1_YN1_MU_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_037:sink_data
	wire          ch1_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                 // id_router_037:sink_ready -> CH1_YN1_MU_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          ch1_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                           // CH1_YN1_ML_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_038:sink_endofpacket
	wire          ch1_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                 // CH1_YN1_ML_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_038:sink_valid
	wire          ch1_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                         // CH1_YN1_ML_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_038:sink_startofpacket
	wire  [102:0] ch1_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rp_data;                                  // CH1_YN1_ML_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_038:sink_data
	wire          ch1_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                 // id_router_038:sink_ready -> CH1_YN1_ML_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          ch1_yn1_l_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                            // CH1_YN1_L_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_039:sink_endofpacket
	wire          ch1_yn1_l_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                  // CH1_YN1_L_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_039:sink_valid
	wire          ch1_yn1_l_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                          // CH1_YN1_L_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_039:sink_startofpacket
	wire  [102:0] ch1_yn1_l_s1_translator_avalon_universal_slave_0_agent_rp_data;                                   // CH1_YN1_L_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_039:sink_data
	wire          ch1_yn1_l_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                  // id_router_039:sink_ready -> CH1_YN1_L_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          ch1_yn2_u_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                            // CH1_YN2_U_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_040:sink_endofpacket
	wire          ch1_yn2_u_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                  // CH1_YN2_U_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_040:sink_valid
	wire          ch1_yn2_u_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                          // CH1_YN2_U_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_040:sink_startofpacket
	wire  [102:0] ch1_yn2_u_s1_translator_avalon_universal_slave_0_agent_rp_data;                                   // CH1_YN2_U_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_040:sink_data
	wire          ch1_yn2_u_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                  // id_router_040:sink_ready -> CH1_YN2_U_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          ch1_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                           // CH1_YN2_MU_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_041:sink_endofpacket
	wire          ch1_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                 // CH1_YN2_MU_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_041:sink_valid
	wire          ch1_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                         // CH1_YN2_MU_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_041:sink_startofpacket
	wire  [102:0] ch1_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rp_data;                                  // CH1_YN2_MU_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_041:sink_data
	wire          ch1_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                 // id_router_041:sink_ready -> CH1_YN2_MU_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          ch1_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                           // CH1_YN2_ML_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_042:sink_endofpacket
	wire          ch1_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                 // CH1_YN2_ML_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_042:sink_valid
	wire          ch1_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                         // CH1_YN2_ML_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_042:sink_startofpacket
	wire  [102:0] ch1_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rp_data;                                  // CH1_YN2_ML_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_042:sink_data
	wire          ch1_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                 // id_router_042:sink_ready -> CH1_YN2_ML_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          ch1_yn2_l_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                            // CH1_YN2_L_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_043:sink_endofpacket
	wire          ch1_yn2_l_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                  // CH1_YN2_L_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_043:sink_valid
	wire          ch1_yn2_l_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                          // CH1_YN2_L_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_043:sink_startofpacket
	wire  [102:0] ch1_yn2_l_s1_translator_avalon_universal_slave_0_agent_rp_data;                                   // CH1_YN2_L_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_043:sink_data
	wire          ch1_yn2_l_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                  // id_router_043:sink_ready -> CH1_YN2_L_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          ch1_yn3_u_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                            // CH1_YN3_U_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_044:sink_endofpacket
	wire          ch1_yn3_u_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                  // CH1_YN3_U_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_044:sink_valid
	wire          ch1_yn3_u_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                          // CH1_YN3_U_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_044:sink_startofpacket
	wire  [102:0] ch1_yn3_u_s1_translator_avalon_universal_slave_0_agent_rp_data;                                   // CH1_YN3_U_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_044:sink_data
	wire          ch1_yn3_u_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                  // id_router_044:sink_ready -> CH1_YN3_U_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          ch1_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                           // CH1_YN3_MU_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_045:sink_endofpacket
	wire          ch1_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                 // CH1_YN3_MU_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_045:sink_valid
	wire          ch1_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                         // CH1_YN3_MU_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_045:sink_startofpacket
	wire  [102:0] ch1_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rp_data;                                  // CH1_YN3_MU_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_045:sink_data
	wire          ch1_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                 // id_router_045:sink_ready -> CH1_YN3_MU_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          ch1_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                           // CH1_YN3_ML_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_046:sink_endofpacket
	wire          ch1_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                 // CH1_YN3_ML_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_046:sink_valid
	wire          ch1_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                         // CH1_YN3_ML_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_046:sink_startofpacket
	wire  [102:0] ch1_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rp_data;                                  // CH1_YN3_ML_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_046:sink_data
	wire          ch1_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                 // id_router_046:sink_ready -> CH1_YN3_ML_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          ch1_yn3_l_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                            // CH1_YN3_L_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_047:sink_endofpacket
	wire          ch1_yn3_l_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                  // CH1_YN3_L_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_047:sink_valid
	wire          ch1_yn3_l_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                          // CH1_YN3_L_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_047:sink_startofpacket
	wire  [102:0] ch1_yn3_l_s1_translator_avalon_universal_slave_0_agent_rp_data;                                   // CH1_YN3_L_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_047:sink_data
	wire          ch1_yn3_l_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                  // id_router_047:sink_ready -> CH1_YN3_L_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          ch2_timer_rst_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                        // CH2_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_048:sink_endofpacket
	wire          ch2_timer_rst_s1_translator_avalon_universal_slave_0_agent_rp_valid;                              // CH2_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_048:sink_valid
	wire          ch2_timer_rst_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                      // CH2_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_048:sink_startofpacket
	wire  [102:0] ch2_timer_rst_s1_translator_avalon_universal_slave_0_agent_rp_data;                               // CH2_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_048:sink_data
	wire          ch2_timer_rst_s1_translator_avalon_universal_slave_0_agent_rp_ready;                              // id_router_048:sink_ready -> CH2_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          ch2_thresh_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                           // CH2_THRESH_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_049:sink_endofpacket
	wire          ch2_thresh_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                 // CH2_THRESH_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_049:sink_valid
	wire          ch2_thresh_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                         // CH2_THRESH_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_049:sink_startofpacket
	wire  [102:0] ch2_thresh_s1_translator_avalon_universal_slave_0_agent_rp_data;                                  // CH2_THRESH_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_049:sink_data
	wire          ch2_thresh_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                 // id_router_049:sink_ready -> CH2_THRESH_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          ch2_rd_peak_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                          // CH2_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_050:sink_endofpacket
	wire          ch2_rd_peak_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                // CH2_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_050:sink_valid
	wire          ch2_rd_peak_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                        // CH2_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_050:sink_startofpacket
	wire  [102:0] ch2_rd_peak_s1_translator_avalon_universal_slave_0_agent_rp_data;                                 // CH2_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_050:sink_data
	wire          ch2_rd_peak_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                // id_router_050:sink_ready -> CH2_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          ch2_peak_found_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                       // CH2_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_051:sink_endofpacket
	wire          ch2_peak_found_s1_translator_avalon_universal_slave_0_agent_rp_valid;                             // CH2_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_051:sink_valid
	wire          ch2_peak_found_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                     // CH2_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_051:sink_startofpacket
	wire  [102:0] ch2_peak_found_s1_translator_avalon_universal_slave_0_agent_rp_data;                              // CH2_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_051:sink_data
	wire          ch2_peak_found_s1_translator_avalon_universal_slave_0_agent_rp_ready;                             // id_router_051:sink_ready -> CH2_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          ch2_time_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                             // CH2_TIME_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_052:sink_endofpacket
	wire          ch2_time_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                   // CH2_TIME_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_052:sink_valid
	wire          ch2_time_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                           // CH2_TIME_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_052:sink_startofpacket
	wire  [102:0] ch2_time_s1_translator_avalon_universal_slave_0_agent_rp_data;                                    // CH2_TIME_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_052:sink_data
	wire          ch2_time_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                   // id_router_052:sink_ready -> CH2_TIME_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          ch2_yn1_u_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                            // CH2_YN1_U_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_053:sink_endofpacket
	wire          ch2_yn1_u_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                  // CH2_YN1_U_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_053:sink_valid
	wire          ch2_yn1_u_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                          // CH2_YN1_U_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_053:sink_startofpacket
	wire  [102:0] ch2_yn1_u_s1_translator_avalon_universal_slave_0_agent_rp_data;                                   // CH2_YN1_U_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_053:sink_data
	wire          ch2_yn1_u_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                  // id_router_053:sink_ready -> CH2_YN1_U_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          ch2_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                           // CH2_YN1_MU_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_054:sink_endofpacket
	wire          ch2_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                 // CH2_YN1_MU_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_054:sink_valid
	wire          ch2_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                         // CH2_YN1_MU_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_054:sink_startofpacket
	wire  [102:0] ch2_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rp_data;                                  // CH2_YN1_MU_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_054:sink_data
	wire          ch2_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                 // id_router_054:sink_ready -> CH2_YN1_MU_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          ch2_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                           // CH2_YN1_ML_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_055:sink_endofpacket
	wire          ch2_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                 // CH2_YN1_ML_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_055:sink_valid
	wire          ch2_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                         // CH2_YN1_ML_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_055:sink_startofpacket
	wire  [102:0] ch2_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rp_data;                                  // CH2_YN1_ML_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_055:sink_data
	wire          ch2_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                 // id_router_055:sink_ready -> CH2_YN1_ML_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          ch2_yn1_l_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                            // CH2_YN1_L_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_056:sink_endofpacket
	wire          ch2_yn1_l_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                  // CH2_YN1_L_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_056:sink_valid
	wire          ch2_yn1_l_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                          // CH2_YN1_L_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_056:sink_startofpacket
	wire  [102:0] ch2_yn1_l_s1_translator_avalon_universal_slave_0_agent_rp_data;                                   // CH2_YN1_L_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_056:sink_data
	wire          ch2_yn1_l_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                  // id_router_056:sink_ready -> CH2_YN1_L_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          ch2_yn2_u_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                            // CH2_YN2_U_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_057:sink_endofpacket
	wire          ch2_yn2_u_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                  // CH2_YN2_U_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_057:sink_valid
	wire          ch2_yn2_u_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                          // CH2_YN2_U_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_057:sink_startofpacket
	wire  [102:0] ch2_yn2_u_s1_translator_avalon_universal_slave_0_agent_rp_data;                                   // CH2_YN2_U_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_057:sink_data
	wire          ch2_yn2_u_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                  // id_router_057:sink_ready -> CH2_YN2_U_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          ch2_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                           // CH2_YN2_MU_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_058:sink_endofpacket
	wire          ch2_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                 // CH2_YN2_MU_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_058:sink_valid
	wire          ch2_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                         // CH2_YN2_MU_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_058:sink_startofpacket
	wire  [102:0] ch2_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rp_data;                                  // CH2_YN2_MU_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_058:sink_data
	wire          ch2_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                 // id_router_058:sink_ready -> CH2_YN2_MU_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          ch2_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                           // CH2_YN2_ML_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_059:sink_endofpacket
	wire          ch2_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                 // CH2_YN2_ML_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_059:sink_valid
	wire          ch2_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                         // CH2_YN2_ML_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_059:sink_startofpacket
	wire  [102:0] ch2_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rp_data;                                  // CH2_YN2_ML_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_059:sink_data
	wire          ch2_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                 // id_router_059:sink_ready -> CH2_YN2_ML_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          ch2_yn2_l_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                            // CH2_YN2_L_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_060:sink_endofpacket
	wire          ch2_yn2_l_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                  // CH2_YN2_L_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_060:sink_valid
	wire          ch2_yn2_l_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                          // CH2_YN2_L_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_060:sink_startofpacket
	wire  [102:0] ch2_yn2_l_s1_translator_avalon_universal_slave_0_agent_rp_data;                                   // CH2_YN2_L_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_060:sink_data
	wire          ch2_yn2_l_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                  // id_router_060:sink_ready -> CH2_YN2_L_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          ch2_yn3_u_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                            // CH2_YN3_U_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_061:sink_endofpacket
	wire          ch2_yn3_u_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                  // CH2_YN3_U_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_061:sink_valid
	wire          ch2_yn3_u_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                          // CH2_YN3_U_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_061:sink_startofpacket
	wire  [102:0] ch2_yn3_u_s1_translator_avalon_universal_slave_0_agent_rp_data;                                   // CH2_YN3_U_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_061:sink_data
	wire          ch2_yn3_u_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                  // id_router_061:sink_ready -> CH2_YN3_U_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          ch2_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                           // CH2_YN3_MU_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_062:sink_endofpacket
	wire          ch2_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                 // CH2_YN3_MU_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_062:sink_valid
	wire          ch2_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                         // CH2_YN3_MU_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_062:sink_startofpacket
	wire  [102:0] ch2_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rp_data;                                  // CH2_YN3_MU_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_062:sink_data
	wire          ch2_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                 // id_router_062:sink_ready -> CH2_YN3_MU_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          ch2_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                           // CH2_YN3_ML_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_063:sink_endofpacket
	wire          ch2_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                 // CH2_YN3_ML_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_063:sink_valid
	wire          ch2_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                         // CH2_YN3_ML_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_063:sink_startofpacket
	wire  [102:0] ch2_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rp_data;                                  // CH2_YN3_ML_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_063:sink_data
	wire          ch2_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                 // id_router_063:sink_ready -> CH2_YN3_ML_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          ch2_yn3_l_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                            // CH2_YN3_L_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_064:sink_endofpacket
	wire          ch2_yn3_l_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                  // CH2_YN3_L_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_064:sink_valid
	wire          ch2_yn3_l_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                          // CH2_YN3_L_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_064:sink_startofpacket
	wire  [102:0] ch2_yn3_l_s1_translator_avalon_universal_slave_0_agent_rp_data;                                   // CH2_YN3_L_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_064:sink_data
	wire          ch2_yn3_l_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                  // id_router_064:sink_ready -> CH2_YN3_L_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          ch3_timer_rst_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                        // CH3_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_065:sink_endofpacket
	wire          ch3_timer_rst_s1_translator_avalon_universal_slave_0_agent_rp_valid;                              // CH3_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_065:sink_valid
	wire          ch3_timer_rst_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                      // CH3_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_065:sink_startofpacket
	wire  [102:0] ch3_timer_rst_s1_translator_avalon_universal_slave_0_agent_rp_data;                               // CH3_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_065:sink_data
	wire          ch3_timer_rst_s1_translator_avalon_universal_slave_0_agent_rp_ready;                              // id_router_065:sink_ready -> CH3_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          ch3_thresh_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                           // CH3_THRESH_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_066:sink_endofpacket
	wire          ch3_thresh_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                 // CH3_THRESH_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_066:sink_valid
	wire          ch3_thresh_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                         // CH3_THRESH_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_066:sink_startofpacket
	wire  [102:0] ch3_thresh_s1_translator_avalon_universal_slave_0_agent_rp_data;                                  // CH3_THRESH_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_066:sink_data
	wire          ch3_thresh_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                 // id_router_066:sink_ready -> CH3_THRESH_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          ch3_rd_peak_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                          // CH3_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_067:sink_endofpacket
	wire          ch3_rd_peak_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                // CH3_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_067:sink_valid
	wire          ch3_rd_peak_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                        // CH3_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_067:sink_startofpacket
	wire  [102:0] ch3_rd_peak_s1_translator_avalon_universal_slave_0_agent_rp_data;                                 // CH3_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_067:sink_data
	wire          ch3_rd_peak_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                // id_router_067:sink_ready -> CH3_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          ch3_peak_found_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                       // CH3_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_068:sink_endofpacket
	wire          ch3_peak_found_s1_translator_avalon_universal_slave_0_agent_rp_valid;                             // CH3_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_068:sink_valid
	wire          ch3_peak_found_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                     // CH3_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_068:sink_startofpacket
	wire  [102:0] ch3_peak_found_s1_translator_avalon_universal_slave_0_agent_rp_data;                              // CH3_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_068:sink_data
	wire          ch3_peak_found_s1_translator_avalon_universal_slave_0_agent_rp_ready;                             // id_router_068:sink_ready -> CH3_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          ch3_yn1_u_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                            // CH3_YN1_U_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_069:sink_endofpacket
	wire          ch3_yn1_u_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                  // CH3_YN1_U_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_069:sink_valid
	wire          ch3_yn1_u_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                          // CH3_YN1_U_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_069:sink_startofpacket
	wire  [102:0] ch3_yn1_u_s1_translator_avalon_universal_slave_0_agent_rp_data;                                   // CH3_YN1_U_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_069:sink_data
	wire          ch3_yn1_u_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                  // id_router_069:sink_ready -> CH3_YN1_U_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          ch3_time_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                             // CH3_TIME_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_070:sink_endofpacket
	wire          ch3_time_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                   // CH3_TIME_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_070:sink_valid
	wire          ch3_time_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                           // CH3_TIME_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_070:sink_startofpacket
	wire  [102:0] ch3_time_s1_translator_avalon_universal_slave_0_agent_rp_data;                                    // CH3_TIME_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_070:sink_data
	wire          ch3_time_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                   // id_router_070:sink_ready -> CH3_TIME_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          ch3_yn3_l_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                            // CH3_YN3_L_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_071:sink_endofpacket
	wire          ch3_yn3_l_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                  // CH3_YN3_L_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_071:sink_valid
	wire          ch3_yn3_l_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                          // CH3_YN3_L_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_071:sink_startofpacket
	wire  [102:0] ch3_yn3_l_s1_translator_avalon_universal_slave_0_agent_rp_data;                                   // CH3_YN3_L_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_071:sink_data
	wire          ch3_yn3_l_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                  // id_router_071:sink_ready -> CH3_YN3_L_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          ch3_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                           // CH3_YN3_ML_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_072:sink_endofpacket
	wire          ch3_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                 // CH3_YN3_ML_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_072:sink_valid
	wire          ch3_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                         // CH3_YN3_ML_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_072:sink_startofpacket
	wire  [102:0] ch3_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rp_data;                                  // CH3_YN3_ML_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_072:sink_data
	wire          ch3_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                 // id_router_072:sink_ready -> CH3_YN3_ML_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          ch3_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                           // CH3_YN3_MU_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_073:sink_endofpacket
	wire          ch3_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                 // CH3_YN3_MU_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_073:sink_valid
	wire          ch3_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                         // CH3_YN3_MU_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_073:sink_startofpacket
	wire  [102:0] ch3_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rp_data;                                  // CH3_YN3_MU_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_073:sink_data
	wire          ch3_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                 // id_router_073:sink_ready -> CH3_YN3_MU_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          ch3_yn3_u_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                            // CH3_YN3_U_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_074:sink_endofpacket
	wire          ch3_yn3_u_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                  // CH3_YN3_U_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_074:sink_valid
	wire          ch3_yn3_u_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                          // CH3_YN3_U_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_074:sink_startofpacket
	wire  [102:0] ch3_yn3_u_s1_translator_avalon_universal_slave_0_agent_rp_data;                                   // CH3_YN3_U_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_074:sink_data
	wire          ch3_yn3_u_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                  // id_router_074:sink_ready -> CH3_YN3_U_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          ch3_yn2_l_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                            // CH3_YN2_L_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_075:sink_endofpacket
	wire          ch3_yn2_l_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                  // CH3_YN2_L_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_075:sink_valid
	wire          ch3_yn2_l_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                          // CH3_YN2_L_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_075:sink_startofpacket
	wire  [102:0] ch3_yn2_l_s1_translator_avalon_universal_slave_0_agent_rp_data;                                   // CH3_YN2_L_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_075:sink_data
	wire          ch3_yn2_l_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                  // id_router_075:sink_ready -> CH3_YN2_L_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          ch3_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                           // CH3_YN2_ML_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_076:sink_endofpacket
	wire          ch3_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                 // CH3_YN2_ML_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_076:sink_valid
	wire          ch3_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                         // CH3_YN2_ML_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_076:sink_startofpacket
	wire  [102:0] ch3_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rp_data;                                  // CH3_YN2_ML_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_076:sink_data
	wire          ch3_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                 // id_router_076:sink_ready -> CH3_YN2_ML_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          ch3_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                           // CH3_YN2_MU_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_077:sink_endofpacket
	wire          ch3_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                 // CH3_YN2_MU_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_077:sink_valid
	wire          ch3_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                         // CH3_YN2_MU_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_077:sink_startofpacket
	wire  [102:0] ch3_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rp_data;                                  // CH3_YN2_MU_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_077:sink_data
	wire          ch3_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                 // id_router_077:sink_ready -> CH3_YN2_MU_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          ch3_yn2_u_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                            // CH3_YN2_U_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_078:sink_endofpacket
	wire          ch3_yn2_u_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                  // CH3_YN2_U_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_078:sink_valid
	wire          ch3_yn2_u_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                          // CH3_YN2_U_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_078:sink_startofpacket
	wire  [102:0] ch3_yn2_u_s1_translator_avalon_universal_slave_0_agent_rp_data;                                   // CH3_YN2_U_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_078:sink_data
	wire          ch3_yn2_u_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                  // id_router_078:sink_ready -> CH3_YN2_U_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          ch3_yn1_l_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                            // CH3_YN1_L_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_079:sink_endofpacket
	wire          ch3_yn1_l_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                  // CH3_YN1_L_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_079:sink_valid
	wire          ch3_yn1_l_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                          // CH3_YN1_L_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_079:sink_startofpacket
	wire  [102:0] ch3_yn1_l_s1_translator_avalon_universal_slave_0_agent_rp_data;                                   // CH3_YN1_L_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_079:sink_data
	wire          ch3_yn1_l_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                  // id_router_079:sink_ready -> CH3_YN1_L_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          ch3_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                           // CH3_YN1_MU_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_080:sink_endofpacket
	wire          ch3_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                 // CH3_YN1_MU_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_080:sink_valid
	wire          ch3_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                         // CH3_YN1_MU_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_080:sink_startofpacket
	wire  [102:0] ch3_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rp_data;                                  // CH3_YN1_MU_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_080:sink_data
	wire          ch3_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                 // id_router_080:sink_ready -> CH3_YN1_MU_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          ch3_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                           // CH3_YN1_ML_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_081:sink_endofpacket
	wire          ch3_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                 // CH3_YN1_ML_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_081:sink_valid
	wire          ch3_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                         // CH3_YN1_ML_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_081:sink_startofpacket
	wire  [102:0] ch3_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rp_data;                                  // CH3_YN1_ML_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_081:sink_data
	wire          ch3_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                 // id_router_081:sink_ready -> CH3_YN1_ML_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          ch4_timer_rst_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                        // CH4_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_082:sink_endofpacket
	wire          ch4_timer_rst_s1_translator_avalon_universal_slave_0_agent_rp_valid;                              // CH4_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_082:sink_valid
	wire          ch4_timer_rst_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                      // CH4_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_082:sink_startofpacket
	wire  [102:0] ch4_timer_rst_s1_translator_avalon_universal_slave_0_agent_rp_data;                               // CH4_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_082:sink_data
	wire          ch4_timer_rst_s1_translator_avalon_universal_slave_0_agent_rp_ready;                              // id_router_082:sink_ready -> CH4_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          ch4_thresh_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                           // CH4_THRESH_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_083:sink_endofpacket
	wire          ch4_thresh_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                 // CH4_THRESH_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_083:sink_valid
	wire          ch4_thresh_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                         // CH4_THRESH_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_083:sink_startofpacket
	wire  [102:0] ch4_thresh_s1_translator_avalon_universal_slave_0_agent_rp_data;                                  // CH4_THRESH_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_083:sink_data
	wire          ch4_thresh_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                 // id_router_083:sink_ready -> CH4_THRESH_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          ch4_rd_peak_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                          // CH4_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_084:sink_endofpacket
	wire          ch4_rd_peak_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                // CH4_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_084:sink_valid
	wire          ch4_rd_peak_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                        // CH4_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_084:sink_startofpacket
	wire  [102:0] ch4_rd_peak_s1_translator_avalon_universal_slave_0_agent_rp_data;                                 // CH4_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_084:sink_data
	wire          ch4_rd_peak_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                // id_router_084:sink_ready -> CH4_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          ch4_peak_found_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                       // CH4_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_085:sink_endofpacket
	wire          ch4_peak_found_s1_translator_avalon_universal_slave_0_agent_rp_valid;                             // CH4_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_085:sink_valid
	wire          ch4_peak_found_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                     // CH4_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_085:sink_startofpacket
	wire  [102:0] ch4_peak_found_s1_translator_avalon_universal_slave_0_agent_rp_data;                              // CH4_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_085:sink_data
	wire          ch4_peak_found_s1_translator_avalon_universal_slave_0_agent_rp_ready;                             // id_router_085:sink_ready -> CH4_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          ch4_time_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                             // CH4_TIME_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_086:sink_endofpacket
	wire          ch4_time_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                   // CH4_TIME_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_086:sink_valid
	wire          ch4_time_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                           // CH4_TIME_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_086:sink_startofpacket
	wire  [102:0] ch4_time_s1_translator_avalon_universal_slave_0_agent_rp_data;                                    // CH4_TIME_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_086:sink_data
	wire          ch4_time_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                   // id_router_086:sink_ready -> CH4_TIME_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          ch4_yn1_u_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                            // CH4_YN1_U_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_087:sink_endofpacket
	wire          ch4_yn1_u_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                  // CH4_YN1_U_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_087:sink_valid
	wire          ch4_yn1_u_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                          // CH4_YN1_U_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_087:sink_startofpacket
	wire  [102:0] ch4_yn1_u_s1_translator_avalon_universal_slave_0_agent_rp_data;                                   // CH4_YN1_U_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_087:sink_data
	wire          ch4_yn1_u_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                  // id_router_087:sink_ready -> CH4_YN1_U_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          ch4_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                           // CH4_YN1_MU_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_088:sink_endofpacket
	wire          ch4_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                 // CH4_YN1_MU_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_088:sink_valid
	wire          ch4_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                         // CH4_YN1_MU_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_088:sink_startofpacket
	wire  [102:0] ch4_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rp_data;                                  // CH4_YN1_MU_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_088:sink_data
	wire          ch4_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                 // id_router_088:sink_ready -> CH4_YN1_MU_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          ch4_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                           // CH4_YN1_ML_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_089:sink_endofpacket
	wire          ch4_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                 // CH4_YN1_ML_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_089:sink_valid
	wire          ch4_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                         // CH4_YN1_ML_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_089:sink_startofpacket
	wire  [102:0] ch4_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rp_data;                                  // CH4_YN1_ML_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_089:sink_data
	wire          ch4_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                 // id_router_089:sink_ready -> CH4_YN1_ML_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          ch4_yn1_l_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                            // CH4_YN1_L_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_090:sink_endofpacket
	wire          ch4_yn1_l_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                  // CH4_YN1_L_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_090:sink_valid
	wire          ch4_yn1_l_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                          // CH4_YN1_L_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_090:sink_startofpacket
	wire  [102:0] ch4_yn1_l_s1_translator_avalon_universal_slave_0_agent_rp_data;                                   // CH4_YN1_L_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_090:sink_data
	wire          ch4_yn1_l_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                  // id_router_090:sink_ready -> CH4_YN1_L_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          ch4_yn2_u_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                            // CH4_YN2_U_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_091:sink_endofpacket
	wire          ch4_yn2_u_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                  // CH4_YN2_U_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_091:sink_valid
	wire          ch4_yn2_u_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                          // CH4_YN2_U_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_091:sink_startofpacket
	wire  [102:0] ch4_yn2_u_s1_translator_avalon_universal_slave_0_agent_rp_data;                                   // CH4_YN2_U_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_091:sink_data
	wire          ch4_yn2_u_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                  // id_router_091:sink_ready -> CH4_YN2_U_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          ch4_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                           // CH4_YN2_MU_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_092:sink_endofpacket
	wire          ch4_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                 // CH4_YN2_MU_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_092:sink_valid
	wire          ch4_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                         // CH4_YN2_MU_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_092:sink_startofpacket
	wire  [102:0] ch4_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rp_data;                                  // CH4_YN2_MU_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_092:sink_data
	wire          ch4_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                 // id_router_092:sink_ready -> CH4_YN2_MU_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          ch4_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                           // CH4_YN2_ML_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_093:sink_endofpacket
	wire          ch4_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                 // CH4_YN2_ML_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_093:sink_valid
	wire          ch4_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                         // CH4_YN2_ML_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_093:sink_startofpacket
	wire  [102:0] ch4_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rp_data;                                  // CH4_YN2_ML_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_093:sink_data
	wire          ch4_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                 // id_router_093:sink_ready -> CH4_YN2_ML_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          ch4_yn2_l_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                            // CH4_YN2_L_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_094:sink_endofpacket
	wire          ch4_yn2_l_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                  // CH4_YN2_L_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_094:sink_valid
	wire          ch4_yn2_l_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                          // CH4_YN2_L_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_094:sink_startofpacket
	wire  [102:0] ch4_yn2_l_s1_translator_avalon_universal_slave_0_agent_rp_data;                                   // CH4_YN2_L_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_094:sink_data
	wire          ch4_yn2_l_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                  // id_router_094:sink_ready -> CH4_YN2_L_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          ch4_yn3_u_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                            // CH4_YN3_U_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_095:sink_endofpacket
	wire          ch4_yn3_u_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                  // CH4_YN3_U_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_095:sink_valid
	wire          ch4_yn3_u_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                          // CH4_YN3_U_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_095:sink_startofpacket
	wire  [102:0] ch4_yn3_u_s1_translator_avalon_universal_slave_0_agent_rp_data;                                   // CH4_YN3_U_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_095:sink_data
	wire          ch4_yn3_u_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                  // id_router_095:sink_ready -> CH4_YN3_U_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          ch4_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                           // CH4_YN3_MU_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_096:sink_endofpacket
	wire          ch4_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                 // CH4_YN3_MU_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_096:sink_valid
	wire          ch4_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                         // CH4_YN3_MU_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_096:sink_startofpacket
	wire  [102:0] ch4_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rp_data;                                  // CH4_YN3_MU_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_096:sink_data
	wire          ch4_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                 // id_router_096:sink_ready -> CH4_YN3_MU_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          ch4_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                           // CH4_YN3_ML_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_097:sink_endofpacket
	wire          ch4_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                 // CH4_YN3_ML_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_097:sink_valid
	wire          ch4_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                         // CH4_YN3_ML_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_097:sink_startofpacket
	wire  [102:0] ch4_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rp_data;                                  // CH4_YN3_ML_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_097:sink_data
	wire          ch4_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                 // id_router_097:sink_ready -> CH4_YN3_ML_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          ch4_yn3_l_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                            // CH4_YN3_L_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_098:sink_endofpacket
	wire          ch4_yn3_l_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                  // CH4_YN3_L_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_098:sink_valid
	wire          ch4_yn3_l_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                          // CH4_YN3_L_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_098:sink_startofpacket
	wire  [102:0] ch4_yn3_l_s1_translator_avalon_universal_slave_0_agent_rp_data;                                   // CH4_YN3_L_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_098:sink_data
	wire          ch4_yn3_l_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                  // id_router_098:sink_ready -> CH4_YN3_L_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          rst_controller_reset_out_reset;                                                                   // rst_controller:reset_out -> [NIOS_CPU:reset_n, NIOS_CPU_data_master_translator:reset, NIOS_CPU_data_master_translator_avalon_universal_master_0_agent:reset, NIOS_CPU_instruction_master_translator:reset, NIOS_CPU_instruction_master_translator_avalon_universal_master_0_agent:reset, NIOS_CPU_jtag_debug_module_translator:reset, NIOS_CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:reset, NIOS_CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, addr_router:reset, addr_router_001:reset, cmd_xbar_demux:reset, cmd_xbar_demux_001:reset, cmd_xbar_mux:reset, id_router:reset, irq_mapper:reset, rsp_xbar_demux:reset, rsp_xbar_mux:reset, rsp_xbar_mux_001:reset]
	wire          rst_controller_001_reset_out_reset;                                                               // rst_controller_001:reset_out -> [ADC_ON:reset_n, ADC_ON_s1_translator:reset, ADC_ON_s1_translator_avalon_universal_slave_0_agent:reset, ADC_ON_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, CH0_PEAK_FOUND:reset_n, CH0_PEAK_FOUND_s1_translator:reset, CH0_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:reset, CH0_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, CH0_RD_PEAK:reset_n, CH0_RD_PEAK_s1_translator:reset, CH0_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:reset, CH0_RD_PEAK_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, CH0_THRESH:reset_n, CH0_THRESH_s1_translator:reset, CH0_THRESH_s1_translator_avalon_universal_slave_0_agent:reset, CH0_THRESH_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, CH0_TIME:reset_n, CH0_TIMER_RST:reset_n, CH0_TIMER_RST_s1_translator:reset, CH0_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:reset, CH0_TIMER_RST_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, CH0_TIME_s1_translator:reset, CH0_TIME_s1_translator_avalon_universal_slave_0_agent:reset, CH0_TIME_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, CH0_YN1_L:reset_n, CH0_YN1_L_s1_translator:reset, CH0_YN1_L_s1_translator_avalon_universal_slave_0_agent:reset, CH0_YN1_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, CH0_YN1_ML:reset_n, CH0_YN1_ML_s1_translator:reset, CH0_YN1_ML_s1_translator_avalon_universal_slave_0_agent:reset, CH0_YN1_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, CH0_YN1_MU:reset_n, CH0_YN1_MU_s1_translator:reset, CH0_YN1_MU_s1_translator_avalon_universal_slave_0_agent:reset, CH0_YN1_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, CH0_YN1_U:reset_n, CH0_YN1_U_s1_translator:reset, CH0_YN1_U_s1_translator_avalon_universal_slave_0_agent:reset, CH0_YN1_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, CH0_YN2_L:reset_n, CH0_YN2_L_s1_translator:reset, CH0_YN2_L_s1_translator_avalon_universal_slave_0_agent:reset, CH0_YN2_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, CH0_YN2_ML:reset_n, CH0_YN2_ML_s1_translator:reset, CH0_YN2_ML_s1_translator_avalon_universal_slave_0_agent:reset, CH0_YN2_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, CH0_YN2_MU:reset_n, CH0_YN2_MU_s1_translator:reset, CH0_YN2_MU_s1_translator_avalon_universal_slave_0_agent:reset, CH0_YN2_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, CH0_YN2_U:reset_n, CH0_YN2_U_s1_translator:reset, CH0_YN2_U_s1_translator_avalon_universal_slave_0_agent:reset, CH0_YN2_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, CH0_YN3_L:reset_n, CH0_YN3_L_s1_translator:reset, CH0_YN3_L_s1_translator_avalon_universal_slave_0_agent:reset, CH0_YN3_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, CH0_YN3_ML:reset_n, CH0_YN3_ML_s1_translator:reset, CH0_YN3_ML_s1_translator_avalon_universal_slave_0_agent:reset, CH0_YN3_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, CH0_YN3_MU:reset_n, CH0_YN3_MU_s1_translator:reset, CH0_YN3_MU_s1_translator_avalon_universal_slave_0_agent:reset, CH0_YN3_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, CH0_YN3_U:reset_n, CH0_YN3_U_s1_translator:reset, CH0_YN3_U_s1_translator_avalon_universal_slave_0_agent:reset, CH0_YN3_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, CH1_PEAK_FOUND:reset_n, CH1_PEAK_FOUND_s1_translator:reset, CH1_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:reset, CH1_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, CH1_RD_PEAK:reset_n, CH1_RD_PEAK_s1_translator:reset, CH1_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:reset, CH1_RD_PEAK_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, CH1_THRESH:reset_n, CH1_THRESH_s1_translator:reset, CH1_THRESH_s1_translator_avalon_universal_slave_0_agent:reset, CH1_THRESH_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, CH1_TIME:reset_n, CH1_TIMER_RST:reset_n, CH1_TIMER_RST_s1_translator:reset, CH1_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:reset, CH1_TIMER_RST_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, CH1_TIME_s1_translator:reset, CH1_TIME_s1_translator_avalon_universal_slave_0_agent:reset, CH1_TIME_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, CH1_YN1_L:reset_n, CH1_YN1_L_s1_translator:reset, CH1_YN1_L_s1_translator_avalon_universal_slave_0_agent:reset, CH1_YN1_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, CH1_YN1_ML:reset_n, CH1_YN1_ML_s1_translator:reset, CH1_YN1_ML_s1_translator_avalon_universal_slave_0_agent:reset, CH1_YN1_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, CH1_YN1_MU:reset_n, CH1_YN1_MU_s1_translator:reset, CH1_YN1_MU_s1_translator_avalon_universal_slave_0_agent:reset, CH1_YN1_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, CH1_YN1_U:reset_n, CH1_YN1_U_s1_translator:reset, CH1_YN1_U_s1_translator_avalon_universal_slave_0_agent:reset, CH1_YN1_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, CH1_YN2_L:reset_n, CH1_YN2_L_s1_translator:reset, CH1_YN2_L_s1_translator_avalon_universal_slave_0_agent:reset, CH1_YN2_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, CH1_YN2_ML:reset_n, CH1_YN2_ML_s1_translator:reset, CH1_YN2_ML_s1_translator_avalon_universal_slave_0_agent:reset, CH1_YN2_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, CH1_YN2_MU:reset_n, CH1_YN2_MU_s1_translator:reset, CH1_YN2_MU_s1_translator_avalon_universal_slave_0_agent:reset, CH1_YN2_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, CH1_YN2_U:reset_n, CH1_YN2_U_s1_translator:reset, CH1_YN2_U_s1_translator_avalon_universal_slave_0_agent:reset, CH1_YN2_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, CH1_YN3_L:reset_n, CH1_YN3_L_s1_translator:reset, CH1_YN3_L_s1_translator_avalon_universal_slave_0_agent:reset, CH1_YN3_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, CH1_YN3_ML:reset_n, CH1_YN3_ML_s1_translator:reset, CH1_YN3_ML_s1_translator_avalon_universal_slave_0_agent:reset, CH1_YN3_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, CH1_YN3_MU:reset_n, CH1_YN3_MU_s1_translator:reset, CH1_YN3_MU_s1_translator_avalon_universal_slave_0_agent:reset, CH1_YN3_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, CH1_YN3_U:reset_n, CH1_YN3_U_s1_translator:reset, CH1_YN3_U_s1_translator_avalon_universal_slave_0_agent:reset, CH1_YN3_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, CH2_PEAK_FOUND:reset_n, CH2_PEAK_FOUND_s1_translator:reset, CH2_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:reset, CH2_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, CH2_RD_PEAK:reset_n, CH2_RD_PEAK_s1_translator:reset, CH2_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:reset, CH2_RD_PEAK_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, CH2_THRESH:reset_n, CH2_THRESH_s1_translator:reset, CH2_THRESH_s1_translator_avalon_universal_slave_0_agent:reset, CH2_THRESH_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, CH2_TIME:reset_n, CH2_TIMER_RST:reset_n, CH2_TIMER_RST_s1_translator:reset, CH2_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:reset, CH2_TIMER_RST_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, CH2_TIME_s1_translator:reset, CH2_TIME_s1_translator_avalon_universal_slave_0_agent:reset, CH2_TIME_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, CH2_YN1_ML:reset_n, CH2_YN1_ML_s1_translator:reset, CH2_YN1_ML_s1_translator_avalon_universal_slave_0_agent:reset, CH2_YN1_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, CH2_YN1_MU:reset_n, CH2_YN1_MU_s1_translator:reset, CH2_YN1_MU_s1_translator_avalon_universal_slave_0_agent:reset, CH2_YN1_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, CH2_YN1_U:reset_n, CH2_YN1_U_s1_translator:reset, CH2_YN1_U_s1_translator_avalon_universal_slave_0_agent:reset, CH2_YN1_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, CH2_YN2_L:reset_n, CH2_YN2_L_s1_translator:reset, CH2_YN2_L_s1_translator_avalon_universal_slave_0_agent:reset, CH2_YN2_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, CH2_YN2_ML:reset_n, CH2_YN2_ML_s1_translator:reset, CH2_YN2_ML_s1_translator_avalon_universal_slave_0_agent:reset, CH2_YN2_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, CH2_YN2_MU:reset_n, CH2_YN2_MU_s1_translator:reset, CH2_YN2_MU_s1_translator_avalon_universal_slave_0_agent:reset, CH2_YN2_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, CH2_YN2_U:reset_n, CH2_YN2_U_s1_translator:reset, CH2_YN2_U_s1_translator_avalon_universal_slave_0_agent:reset, CH2_YN2_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, CH2_YN3_L:reset_n, CH2_YN3_L_s1_translator:reset, CH2_YN3_L_s1_translator_avalon_universal_slave_0_agent:reset, CH2_YN3_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, CH2_YN3_ML:reset_n, CH2_YN3_ML_s1_translator:reset, CH2_YN3_ML_s1_translator_avalon_universal_slave_0_agent:reset, CH2_YN3_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, CH2_YN3_MU:reset_n, CH2_YN3_MU_s1_translator:reset, CH2_YN3_MU_s1_translator_avalon_universal_slave_0_agent:reset, CH2_YN3_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, CH2_YN3_U:reset_n, CH2_YN3_U_s1_translator:reset, CH2_YN3_U_s1_translator_avalon_universal_slave_0_agent:reset, CH2_YN3_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, CH3_PEAK_FOUND:reset_n, CH3_PEAK_FOUND_s1_translator:reset, CH3_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:reset, CH3_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, CH3_RD_PEAK:reset_n, CH3_RD_PEAK_s1_translator:reset, CH3_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:reset, CH3_RD_PEAK_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, CH3_THRESH:reset_n, CH3_THRESH_s1_translator:reset, CH3_THRESH_s1_translator_avalon_universal_slave_0_agent:reset, CH3_THRESH_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, CH3_TIME:reset_n, CH3_TIMER_RST:reset_n, CH3_TIMER_RST_s1_translator:reset, CH3_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:reset, CH3_TIMER_RST_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, CH3_TIME_s1_translator:reset, CH3_TIME_s1_translator_avalon_universal_slave_0_agent:reset, CH3_TIME_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, CH3_YN1_L:reset_n, CH3_YN1_L_s1_translator:reset, CH3_YN1_L_s1_translator_avalon_universal_slave_0_agent:reset, CH3_YN1_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, CH3_YN1_ML:reset_n, CH3_YN1_ML_s1_translator:reset, CH3_YN1_ML_s1_translator_avalon_universal_slave_0_agent:reset, CH3_YN1_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, CH3_YN1_MU:reset_n, CH3_YN1_MU_s1_translator:reset, CH3_YN1_MU_s1_translator_avalon_universal_slave_0_agent:reset, CH3_YN1_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, CH3_YN1_U:reset_n, CH3_YN1_U_s1_translator:reset, CH3_YN1_U_s1_translator_avalon_universal_slave_0_agent:reset, CH3_YN1_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, CH3_YN2_L:reset_n, CH3_YN2_L_s1_translator:reset, CH3_YN2_L_s1_translator_avalon_universal_slave_0_agent:reset, CH3_YN2_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, CH3_YN2_ML:reset_n, CH3_YN2_ML_s1_translator:reset, CH3_YN2_ML_s1_translator_avalon_universal_slave_0_agent:reset, CH3_YN2_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, CH3_YN2_MU:reset_n, CH3_YN2_MU_s1_translator:reset, CH3_YN2_MU_s1_translator_avalon_universal_slave_0_agent:reset, CH3_YN2_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, CH3_YN2_U:reset_n, CH3_YN2_U_s1_translator:reset, CH3_YN2_U_s1_translator_avalon_universal_slave_0_agent:reset, CH3_YN2_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, CH3_YN3_L:reset_n, CH3_YN3_L_s1_translator:reset, CH3_YN3_L_s1_translator_avalon_universal_slave_0_agent:reset, CH3_YN3_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, CH3_YN3_ML:reset_n, CH3_YN3_ML_s1_translator:reset, CH3_YN3_ML_s1_translator_avalon_universal_slave_0_agent:reset, CH3_YN3_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, CH3_YN3_MU:reset_n, CH3_YN3_MU_s1_translator:reset, CH3_YN3_MU_s1_translator_avalon_universal_slave_0_agent:reset, CH3_YN3_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, CH3_YN3_U:reset_n, CH3_YN3_U_s1_translator:reset, CH3_YN3_U_s1_translator_avalon_universal_slave_0_agent:reset, CH3_YN3_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, CH4_PEAK_FOUND:reset_n, CH4_PEAK_FOUND_s1_translator:reset, CH4_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:reset, CH4_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, CH4_RD_PEAK:reset_n, CH4_RD_PEAK_s1_translator:reset, CH4_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:reset, CH4_RD_PEAK_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, CH4_THRESH:reset_n, CH4_THRESH_s1_translator:reset, CH4_THRESH_s1_translator_avalon_universal_slave_0_agent:reset, CH4_THRESH_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, CH4_TIME:reset_n, CH4_TIMER_RST:reset_n, CH4_TIMER_RST_s1_translator:reset, CH4_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:reset, CH4_TIMER_RST_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, CH4_TIME_s1_translator:reset, CH4_TIME_s1_translator_avalon_universal_slave_0_agent:reset, CH4_TIME_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, CH4_YN1_L:reset_n, CH4_YN1_L_s1_translator:reset, CH4_YN1_L_s1_translator_avalon_universal_slave_0_agent:reset, CH4_YN1_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, CH4_YN1_ML:reset_n, CH4_YN1_ML_s1_translator:reset, CH4_YN1_ML_s1_translator_avalon_universal_slave_0_agent:reset, CH4_YN1_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, CH4_YN1_MU:reset_n, CH4_YN1_MU_s1_translator:reset, CH4_YN1_MU_s1_translator_avalon_universal_slave_0_agent:reset, CH4_YN1_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, CH4_YN1_U:reset_n, CH4_YN1_U_s1_translator:reset, CH4_YN1_U_s1_translator_avalon_universal_slave_0_agent:reset, CH4_YN1_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, CH4_YN2_L:reset_n, CH4_YN2_L_s1_translator:reset, CH4_YN2_L_s1_translator_avalon_universal_slave_0_agent:reset, CH4_YN2_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, CH4_YN2_ML:reset_n, CH4_YN2_ML_s1_translator:reset, CH4_YN2_ML_s1_translator_avalon_universal_slave_0_agent:reset, CH4_YN2_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, CH4_YN2_MU:reset_n, CH4_YN2_MU_s1_translator:reset, CH4_YN2_MU_s1_translator_avalon_universal_slave_0_agent:reset, CH4_YN2_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, CH4_YN2_U:reset_n, CH4_YN2_U_s1_translator:reset, CH4_YN2_U_s1_translator_avalon_universal_slave_0_agent:reset, CH4_YN2_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, CH4_YN3_L:reset_n, CH4_YN3_L_s1_translator:reset, CH4_YN3_L_s1_translator_avalon_universal_slave_0_agent:reset, CH4_YN3_L_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, CH4_YN3_ML:reset_n, CH4_YN3_ML_s1_translator:reset, CH4_YN3_ML_s1_translator_avalon_universal_slave_0_agent:reset, CH4_YN3_ML_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, CH4_YN3_MU:reset_n, CH4_YN3_MU_s1_translator:reset, CH4_YN3_MU_s1_translator_avalon_universal_slave_0_agent:reset, CH4_YN3_MU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, CH4_YN3_U:reset_n, CH4_YN3_U_s1_translator:reset, CH4_YN3_U_s1_translator_avalon_universal_slave_0_agent:reset, CH4_YN3_U_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, DETECTOR_ON:reset_n, DETECTOR_ON_s1_translator:reset, DETECTOR_ON_s1_translator_avalon_universal_slave_0_agent:reset, DETECTOR_ON_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, FIFO_ADC_DATA:reset_n, FIFO_ADC_DATA_VALID:reset_n, FIFO_ADC_DATA_VALID_s1_translator:reset, FIFO_ADC_DATA_VALID_s1_translator_avalon_universal_slave_0_agent:reset, FIFO_ADC_DATA_VALID_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, FIFO_ADC_DATA_s1_translator:reset, FIFO_ADC_DATA_s1_translator_avalon_universal_slave_0_agent:reset, FIFO_ADC_DATA_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, FIFO_RST:reset_n, FIFO_RST_s1_translator:reset, FIFO_RST_s1_translator_avalon_universal_slave_0_agent:reset, FIFO_RST_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, JTAG_UART:rst_n, JTAG_UART_avalon_jtag_slave_translator:reset, JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:reset, JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, LCD:reset_n, LCD_control_slave_translator:reset, LCD_control_slave_translator_avalon_universal_slave_0_agent:reset, LCD_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, MENU:reset_n, MENU_DOWN:reset_n, MENU_DOWN_s1_translator:reset, MENU_DOWN_s1_translator_avalon_universal_slave_0_agent:reset, MENU_DOWN_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, MENU_UP:reset_n, MENU_UP_s1_translator:reset, MENU_UP_s1_translator_avalon_universal_slave_0_agent:reset, MENU_UP_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, MENU_s1_translator:reset, MENU_s1_translator_avalon_universal_slave_0_agent:reset, MENU_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, RAM:reset, RAM_s1_translator:reset, RAM_s1_translator_avalon_universal_slave_0_agent:reset, RAM_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, SSRAM:reset_reset, SSRAM_uas_translator:reset, SSRAM_uas_translator_avalon_universal_slave_0_agent:reset, SSRAM_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, SUBTRACTOR_ON:reset_n, SUBTRACTOR_ON_s1_translator:reset, SUBTRACTOR_ON_s1_translator_avalon_universal_slave_0_agent:reset, SUBTRACTOR_ON_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, cmd_xbar_mux_001:reset, cmd_xbar_mux_002:reset, id_router_001:reset, id_router_002:reset, id_router_003:reset, id_router_004:reset, id_router_005:reset, id_router_006:reset, id_router_007:reset, id_router_008:reset, id_router_009:reset, id_router_010:reset, id_router_011:reset, id_router_012:reset, id_router_013:reset, id_router_014:reset, id_router_015:reset, id_router_016:reset, id_router_017:reset, id_router_018:reset, id_router_019:reset, id_router_020:reset, id_router_021:reset, id_router_022:reset, id_router_023:reset, id_router_024:reset, id_router_025:reset, id_router_026:reset, id_router_027:reset, id_router_028:reset, id_router_029:reset, id_router_030:reset, id_router_031:reset, id_router_032:reset, id_router_033:reset, id_router_034:reset, id_router_035:reset, id_router_036:reset, id_router_037:reset, id_router_038:reset, id_router_039:reset, id_router_040:reset, id_router_041:reset, id_router_042:reset, id_router_043:reset, id_router_044:reset, id_router_045:reset, id_router_046:reset, id_router_047:reset, id_router_048:reset, id_router_049:reset, id_router_050:reset, id_router_051:reset, id_router_052:reset, id_router_053:reset, id_router_054:reset, id_router_055:reset, id_router_057:reset, id_router_058:reset, id_router_059:reset, id_router_060:reset, id_router_061:reset, id_router_062:reset, id_router_063:reset, id_router_064:reset, id_router_065:reset, id_router_066:reset, id_router_067:reset, id_router_068:reset, id_router_069:reset, id_router_070:reset, id_router_071:reset, id_router_072:reset, id_router_073:reset, id_router_074:reset, id_router_075:reset, id_router_076:reset, id_router_077:reset, id_router_078:reset, id_router_079:reset, id_router_080:reset, id_router_081:reset, id_router_082:reset, id_router_083:reset, id_router_084:reset, id_router_085:reset, id_router_086:reset, id_router_087:reset, id_router_088:reset, id_router_089:reset, id_router_090:reset, id_router_091:reset, id_router_092:reset, id_router_093:reset, id_router_094:reset, id_router_095:reset, id_router_096:reset, id_router_097:reset, id_router_098:reset, rsp_xbar_demux_001:reset, rsp_xbar_demux_002:reset, rsp_xbar_demux_003:reset, rsp_xbar_demux_004:reset, rsp_xbar_demux_005:reset, rsp_xbar_demux_006:reset, rsp_xbar_demux_007:reset, rsp_xbar_demux_008:reset, rsp_xbar_demux_009:reset, rsp_xbar_demux_010:reset, rsp_xbar_demux_011:reset, rsp_xbar_demux_012:reset, rsp_xbar_demux_013:reset, rsp_xbar_demux_014:reset, rsp_xbar_demux_015:reset, rsp_xbar_demux_016:reset, rsp_xbar_demux_017:reset, rsp_xbar_demux_018:reset, rsp_xbar_demux_019:reset, rsp_xbar_demux_020:reset, rsp_xbar_demux_021:reset, rsp_xbar_demux_022:reset, rsp_xbar_demux_023:reset, rsp_xbar_demux_024:reset, rsp_xbar_demux_025:reset, rsp_xbar_demux_026:reset, rsp_xbar_demux_027:reset, rsp_xbar_demux_028:reset, rsp_xbar_demux_029:reset, rsp_xbar_demux_030:reset, rsp_xbar_demux_031:reset, rsp_xbar_demux_032:reset, rsp_xbar_demux_033:reset, rsp_xbar_demux_034:reset, rsp_xbar_demux_035:reset, rsp_xbar_demux_036:reset, rsp_xbar_demux_037:reset, rsp_xbar_demux_038:reset, rsp_xbar_demux_039:reset, rsp_xbar_demux_040:reset, rsp_xbar_demux_041:reset, rsp_xbar_demux_042:reset, rsp_xbar_demux_043:reset, rsp_xbar_demux_044:reset, rsp_xbar_demux_045:reset, rsp_xbar_demux_046:reset, rsp_xbar_demux_047:reset, rsp_xbar_demux_048:reset, rsp_xbar_demux_049:reset, rsp_xbar_demux_050:reset, rsp_xbar_demux_051:reset, rsp_xbar_demux_052:reset, rsp_xbar_demux_053:reset, rsp_xbar_demux_054:reset, rsp_xbar_demux_055:reset, rsp_xbar_demux_057:reset, rsp_xbar_demux_058:reset, rsp_xbar_demux_059:reset, rsp_xbar_demux_060:reset, rsp_xbar_demux_061:reset, rsp_xbar_demux_062:reset, rsp_xbar_demux_063:reset, rsp_xbar_demux_064:reset, rsp_xbar_demux_065:reset, rsp_xbar_demux_066:reset, rsp_xbar_demux_067:reset, rsp_xbar_demux_068:reset, rsp_xbar_demux_069:reset, rsp_xbar_demux_070:reset, rsp_xbar_demux_071:reset, rsp_xbar_demux_072:reset, rsp_xbar_demux_073:reset, rsp_xbar_demux_074:reset, rsp_xbar_demux_075:reset, rsp_xbar_demux_076:reset, rsp_xbar_demux_077:reset, rsp_xbar_demux_078:reset, rsp_xbar_demux_079:reset, rsp_xbar_demux_080:reset, rsp_xbar_demux_081:reset, rsp_xbar_demux_082:reset, rsp_xbar_demux_083:reset, rsp_xbar_demux_084:reset, rsp_xbar_demux_085:reset, rsp_xbar_demux_086:reset, rsp_xbar_demux_087:reset, rsp_xbar_demux_088:reset, rsp_xbar_demux_089:reset, rsp_xbar_demux_090:reset, rsp_xbar_demux_091:reset, rsp_xbar_demux_092:reset, rsp_xbar_demux_093:reset, rsp_xbar_demux_094:reset, rsp_xbar_demux_095:reset, rsp_xbar_demux_096:reset, rsp_xbar_demux_097:reset, rsp_xbar_demux_098:reset, tristate_bridge_ssram:reset, tristate_bridge_ssram_pinSharer:reset_reset]
	wire          rst_controller_001_reset_out_reset_req;                                                           // rst_controller_001:reset_req -> RAM:reset_req
	wire          cmd_xbar_demux_src0_endofpacket;                                                                  // cmd_xbar_demux:src0_endofpacket -> cmd_xbar_mux:sink0_endofpacket
	wire          cmd_xbar_demux_src0_valid;                                                                        // cmd_xbar_demux:src0_valid -> cmd_xbar_mux:sink0_valid
	wire          cmd_xbar_demux_src0_startofpacket;                                                                // cmd_xbar_demux:src0_startofpacket -> cmd_xbar_mux:sink0_startofpacket
	wire  [102:0] cmd_xbar_demux_src0_data;                                                                         // cmd_xbar_demux:src0_data -> cmd_xbar_mux:sink0_data
	wire   [98:0] cmd_xbar_demux_src0_channel;                                                                      // cmd_xbar_demux:src0_channel -> cmd_xbar_mux:sink0_channel
	wire          cmd_xbar_demux_src0_ready;                                                                        // cmd_xbar_mux:sink0_ready -> cmd_xbar_demux:src0_ready
	wire          cmd_xbar_demux_src1_endofpacket;                                                                  // cmd_xbar_demux:src1_endofpacket -> cmd_xbar_mux_001:sink0_endofpacket
	wire          cmd_xbar_demux_src1_valid;                                                                        // cmd_xbar_demux:src1_valid -> cmd_xbar_mux_001:sink0_valid
	wire          cmd_xbar_demux_src1_startofpacket;                                                                // cmd_xbar_demux:src1_startofpacket -> cmd_xbar_mux_001:sink0_startofpacket
	wire  [102:0] cmd_xbar_demux_src1_data;                                                                         // cmd_xbar_demux:src1_data -> cmd_xbar_mux_001:sink0_data
	wire   [98:0] cmd_xbar_demux_src1_channel;                                                                      // cmd_xbar_demux:src1_channel -> cmd_xbar_mux_001:sink0_channel
	wire          cmd_xbar_demux_src1_ready;                                                                        // cmd_xbar_mux_001:sink0_ready -> cmd_xbar_demux:src1_ready
	wire          cmd_xbar_demux_src2_endofpacket;                                                                  // cmd_xbar_demux:src2_endofpacket -> cmd_xbar_mux_002:sink0_endofpacket
	wire          cmd_xbar_demux_src2_valid;                                                                        // cmd_xbar_demux:src2_valid -> cmd_xbar_mux_002:sink0_valid
	wire          cmd_xbar_demux_src2_startofpacket;                                                                // cmd_xbar_demux:src2_startofpacket -> cmd_xbar_mux_002:sink0_startofpacket
	wire  [102:0] cmd_xbar_demux_src2_data;                                                                         // cmd_xbar_demux:src2_data -> cmd_xbar_mux_002:sink0_data
	wire   [98:0] cmd_xbar_demux_src2_channel;                                                                      // cmd_xbar_demux:src2_channel -> cmd_xbar_mux_002:sink0_channel
	wire          cmd_xbar_demux_src2_ready;                                                                        // cmd_xbar_mux_002:sink0_ready -> cmd_xbar_demux:src2_ready
	wire          cmd_xbar_demux_001_src0_endofpacket;                                                              // cmd_xbar_demux_001:src0_endofpacket -> cmd_xbar_mux:sink1_endofpacket
	wire          cmd_xbar_demux_001_src0_valid;                                                                    // cmd_xbar_demux_001:src0_valid -> cmd_xbar_mux:sink1_valid
	wire          cmd_xbar_demux_001_src0_startofpacket;                                                            // cmd_xbar_demux_001:src0_startofpacket -> cmd_xbar_mux:sink1_startofpacket
	wire  [102:0] cmd_xbar_demux_001_src0_data;                                                                     // cmd_xbar_demux_001:src0_data -> cmd_xbar_mux:sink1_data
	wire   [98:0] cmd_xbar_demux_001_src0_channel;                                                                  // cmd_xbar_demux_001:src0_channel -> cmd_xbar_mux:sink1_channel
	wire          cmd_xbar_demux_001_src0_ready;                                                                    // cmd_xbar_mux:sink1_ready -> cmd_xbar_demux_001:src0_ready
	wire          cmd_xbar_demux_001_src1_endofpacket;                                                              // cmd_xbar_demux_001:src1_endofpacket -> cmd_xbar_mux_001:sink1_endofpacket
	wire          cmd_xbar_demux_001_src1_valid;                                                                    // cmd_xbar_demux_001:src1_valid -> cmd_xbar_mux_001:sink1_valid
	wire          cmd_xbar_demux_001_src1_startofpacket;                                                            // cmd_xbar_demux_001:src1_startofpacket -> cmd_xbar_mux_001:sink1_startofpacket
	wire  [102:0] cmd_xbar_demux_001_src1_data;                                                                     // cmd_xbar_demux_001:src1_data -> cmd_xbar_mux_001:sink1_data
	wire   [98:0] cmd_xbar_demux_001_src1_channel;                                                                  // cmd_xbar_demux_001:src1_channel -> cmd_xbar_mux_001:sink1_channel
	wire          cmd_xbar_demux_001_src1_ready;                                                                    // cmd_xbar_mux_001:sink1_ready -> cmd_xbar_demux_001:src1_ready
	wire          cmd_xbar_demux_001_src2_endofpacket;                                                              // cmd_xbar_demux_001:src2_endofpacket -> cmd_xbar_mux_002:sink1_endofpacket
	wire          cmd_xbar_demux_001_src2_valid;                                                                    // cmd_xbar_demux_001:src2_valid -> cmd_xbar_mux_002:sink1_valid
	wire          cmd_xbar_demux_001_src2_startofpacket;                                                            // cmd_xbar_demux_001:src2_startofpacket -> cmd_xbar_mux_002:sink1_startofpacket
	wire  [102:0] cmd_xbar_demux_001_src2_data;                                                                     // cmd_xbar_demux_001:src2_data -> cmd_xbar_mux_002:sink1_data
	wire   [98:0] cmd_xbar_demux_001_src2_channel;                                                                  // cmd_xbar_demux_001:src2_channel -> cmd_xbar_mux_002:sink1_channel
	wire          cmd_xbar_demux_001_src2_ready;                                                                    // cmd_xbar_mux_002:sink1_ready -> cmd_xbar_demux_001:src2_ready
	wire          cmd_xbar_demux_001_src3_endofpacket;                                                              // cmd_xbar_demux_001:src3_endofpacket -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src3_valid;                                                                    // cmd_xbar_demux_001:src3_valid -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src3_startofpacket;                                                            // cmd_xbar_demux_001:src3_startofpacket -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] cmd_xbar_demux_001_src3_data;                                                                     // cmd_xbar_demux_001:src3_data -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [98:0] cmd_xbar_demux_001_src3_channel;                                                                  // cmd_xbar_demux_001:src3_channel -> JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src4_endofpacket;                                                              // cmd_xbar_demux_001:src4_endofpacket -> LCD_control_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src4_valid;                                                                    // cmd_xbar_demux_001:src4_valid -> LCD_control_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src4_startofpacket;                                                            // cmd_xbar_demux_001:src4_startofpacket -> LCD_control_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] cmd_xbar_demux_001_src4_data;                                                                     // cmd_xbar_demux_001:src4_data -> LCD_control_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [98:0] cmd_xbar_demux_001_src4_channel;                                                                  // cmd_xbar_demux_001:src4_channel -> LCD_control_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src5_endofpacket;                                                              // cmd_xbar_demux_001:src5_endofpacket -> ADC_ON_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src5_valid;                                                                    // cmd_xbar_demux_001:src5_valid -> ADC_ON_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src5_startofpacket;                                                            // cmd_xbar_demux_001:src5_startofpacket -> ADC_ON_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] cmd_xbar_demux_001_src5_data;                                                                     // cmd_xbar_demux_001:src5_data -> ADC_ON_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [98:0] cmd_xbar_demux_001_src5_channel;                                                                  // cmd_xbar_demux_001:src5_channel -> ADC_ON_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src6_endofpacket;                                                              // cmd_xbar_demux_001:src6_endofpacket -> FIFO_ADC_DATA_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src6_valid;                                                                    // cmd_xbar_demux_001:src6_valid -> FIFO_ADC_DATA_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src6_startofpacket;                                                            // cmd_xbar_demux_001:src6_startofpacket -> FIFO_ADC_DATA_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] cmd_xbar_demux_001_src6_data;                                                                     // cmd_xbar_demux_001:src6_data -> FIFO_ADC_DATA_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [98:0] cmd_xbar_demux_001_src6_channel;                                                                  // cmd_xbar_demux_001:src6_channel -> FIFO_ADC_DATA_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src7_endofpacket;                                                              // cmd_xbar_demux_001:src7_endofpacket -> FIFO_ADC_DATA_VALID_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src7_valid;                                                                    // cmd_xbar_demux_001:src7_valid -> FIFO_ADC_DATA_VALID_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src7_startofpacket;                                                            // cmd_xbar_demux_001:src7_startofpacket -> FIFO_ADC_DATA_VALID_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] cmd_xbar_demux_001_src7_data;                                                                     // cmd_xbar_demux_001:src7_data -> FIFO_ADC_DATA_VALID_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [98:0] cmd_xbar_demux_001_src7_channel;                                                                  // cmd_xbar_demux_001:src7_channel -> FIFO_ADC_DATA_VALID_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src8_endofpacket;                                                              // cmd_xbar_demux_001:src8_endofpacket -> FIFO_RST_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src8_valid;                                                                    // cmd_xbar_demux_001:src8_valid -> FIFO_RST_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src8_startofpacket;                                                            // cmd_xbar_demux_001:src8_startofpacket -> FIFO_RST_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] cmd_xbar_demux_001_src8_data;                                                                     // cmd_xbar_demux_001:src8_data -> FIFO_RST_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [98:0] cmd_xbar_demux_001_src8_channel;                                                                  // cmd_xbar_demux_001:src8_channel -> FIFO_RST_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src9_endofpacket;                                                              // cmd_xbar_demux_001:src9_endofpacket -> SUBTRACTOR_ON_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src9_valid;                                                                    // cmd_xbar_demux_001:src9_valid -> SUBTRACTOR_ON_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src9_startofpacket;                                                            // cmd_xbar_demux_001:src9_startofpacket -> SUBTRACTOR_ON_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] cmd_xbar_demux_001_src9_data;                                                                     // cmd_xbar_demux_001:src9_data -> SUBTRACTOR_ON_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [98:0] cmd_xbar_demux_001_src9_channel;                                                                  // cmd_xbar_demux_001:src9_channel -> SUBTRACTOR_ON_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src10_endofpacket;                                                             // cmd_xbar_demux_001:src10_endofpacket -> CH0_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src10_valid;                                                                   // cmd_xbar_demux_001:src10_valid -> CH0_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src10_startofpacket;                                                           // cmd_xbar_demux_001:src10_startofpacket -> CH0_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] cmd_xbar_demux_001_src10_data;                                                                    // cmd_xbar_demux_001:src10_data -> CH0_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [98:0] cmd_xbar_demux_001_src10_channel;                                                                 // cmd_xbar_demux_001:src10_channel -> CH0_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src11_endofpacket;                                                             // cmd_xbar_demux_001:src11_endofpacket -> DETECTOR_ON_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src11_valid;                                                                   // cmd_xbar_demux_001:src11_valid -> DETECTOR_ON_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src11_startofpacket;                                                           // cmd_xbar_demux_001:src11_startofpacket -> DETECTOR_ON_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] cmd_xbar_demux_001_src11_data;                                                                    // cmd_xbar_demux_001:src11_data -> DETECTOR_ON_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [98:0] cmd_xbar_demux_001_src11_channel;                                                                 // cmd_xbar_demux_001:src11_channel -> DETECTOR_ON_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src12_endofpacket;                                                             // cmd_xbar_demux_001:src12_endofpacket -> MENU_DOWN_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src12_valid;                                                                   // cmd_xbar_demux_001:src12_valid -> MENU_DOWN_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src12_startofpacket;                                                           // cmd_xbar_demux_001:src12_startofpacket -> MENU_DOWN_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] cmd_xbar_demux_001_src12_data;                                                                    // cmd_xbar_demux_001:src12_data -> MENU_DOWN_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [98:0] cmd_xbar_demux_001_src12_channel;                                                                 // cmd_xbar_demux_001:src12_channel -> MENU_DOWN_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src13_endofpacket;                                                             // cmd_xbar_demux_001:src13_endofpacket -> MENU_UP_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src13_valid;                                                                   // cmd_xbar_demux_001:src13_valid -> MENU_UP_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src13_startofpacket;                                                           // cmd_xbar_demux_001:src13_startofpacket -> MENU_UP_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] cmd_xbar_demux_001_src13_data;                                                                    // cmd_xbar_demux_001:src13_data -> MENU_UP_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [98:0] cmd_xbar_demux_001_src13_channel;                                                                 // cmd_xbar_demux_001:src13_channel -> MENU_UP_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src14_endofpacket;                                                             // cmd_xbar_demux_001:src14_endofpacket -> MENU_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src14_valid;                                                                   // cmd_xbar_demux_001:src14_valid -> MENU_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src14_startofpacket;                                                           // cmd_xbar_demux_001:src14_startofpacket -> MENU_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] cmd_xbar_demux_001_src14_data;                                                                    // cmd_xbar_demux_001:src14_data -> MENU_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [98:0] cmd_xbar_demux_001_src14_channel;                                                                 // cmd_xbar_demux_001:src14_channel -> MENU_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src15_endofpacket;                                                             // cmd_xbar_demux_001:src15_endofpacket -> CH0_THRESH_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src15_valid;                                                                   // cmd_xbar_demux_001:src15_valid -> CH0_THRESH_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src15_startofpacket;                                                           // cmd_xbar_demux_001:src15_startofpacket -> CH0_THRESH_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] cmd_xbar_demux_001_src15_data;                                                                    // cmd_xbar_demux_001:src15_data -> CH0_THRESH_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [98:0] cmd_xbar_demux_001_src15_channel;                                                                 // cmd_xbar_demux_001:src15_channel -> CH0_THRESH_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src16_endofpacket;                                                             // cmd_xbar_demux_001:src16_endofpacket -> CH0_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src16_valid;                                                                   // cmd_xbar_demux_001:src16_valid -> CH0_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src16_startofpacket;                                                           // cmd_xbar_demux_001:src16_startofpacket -> CH0_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] cmd_xbar_demux_001_src16_data;                                                                    // cmd_xbar_demux_001:src16_data -> CH0_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [98:0] cmd_xbar_demux_001_src16_channel;                                                                 // cmd_xbar_demux_001:src16_channel -> CH0_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src17_endofpacket;                                                             // cmd_xbar_demux_001:src17_endofpacket -> CH0_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src17_valid;                                                                   // cmd_xbar_demux_001:src17_valid -> CH0_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src17_startofpacket;                                                           // cmd_xbar_demux_001:src17_startofpacket -> CH0_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] cmd_xbar_demux_001_src17_data;                                                                    // cmd_xbar_demux_001:src17_data -> CH0_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [98:0] cmd_xbar_demux_001_src17_channel;                                                                 // cmd_xbar_demux_001:src17_channel -> CH0_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src18_endofpacket;                                                             // cmd_xbar_demux_001:src18_endofpacket -> CH0_YN1_L_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src18_valid;                                                                   // cmd_xbar_demux_001:src18_valid -> CH0_YN1_L_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src18_startofpacket;                                                           // cmd_xbar_demux_001:src18_startofpacket -> CH0_YN1_L_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] cmd_xbar_demux_001_src18_data;                                                                    // cmd_xbar_demux_001:src18_data -> CH0_YN1_L_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [98:0] cmd_xbar_demux_001_src18_channel;                                                                 // cmd_xbar_demux_001:src18_channel -> CH0_YN1_L_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src19_endofpacket;                                                             // cmd_xbar_demux_001:src19_endofpacket -> CH0_YN1_ML_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src19_valid;                                                                   // cmd_xbar_demux_001:src19_valid -> CH0_YN1_ML_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src19_startofpacket;                                                           // cmd_xbar_demux_001:src19_startofpacket -> CH0_YN1_ML_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] cmd_xbar_demux_001_src19_data;                                                                    // cmd_xbar_demux_001:src19_data -> CH0_YN1_ML_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [98:0] cmd_xbar_demux_001_src19_channel;                                                                 // cmd_xbar_demux_001:src19_channel -> CH0_YN1_ML_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src20_endofpacket;                                                             // cmd_xbar_demux_001:src20_endofpacket -> CH0_YN1_MU_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src20_valid;                                                                   // cmd_xbar_demux_001:src20_valid -> CH0_YN1_MU_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src20_startofpacket;                                                           // cmd_xbar_demux_001:src20_startofpacket -> CH0_YN1_MU_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] cmd_xbar_demux_001_src20_data;                                                                    // cmd_xbar_demux_001:src20_data -> CH0_YN1_MU_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [98:0] cmd_xbar_demux_001_src20_channel;                                                                 // cmd_xbar_demux_001:src20_channel -> CH0_YN1_MU_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src21_endofpacket;                                                             // cmd_xbar_demux_001:src21_endofpacket -> CH0_YN1_U_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src21_valid;                                                                   // cmd_xbar_demux_001:src21_valid -> CH0_YN1_U_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src21_startofpacket;                                                           // cmd_xbar_demux_001:src21_startofpacket -> CH0_YN1_U_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] cmd_xbar_demux_001_src21_data;                                                                    // cmd_xbar_demux_001:src21_data -> CH0_YN1_U_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [98:0] cmd_xbar_demux_001_src21_channel;                                                                 // cmd_xbar_demux_001:src21_channel -> CH0_YN1_U_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src22_endofpacket;                                                             // cmd_xbar_demux_001:src22_endofpacket -> CH0_TIME_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src22_valid;                                                                   // cmd_xbar_demux_001:src22_valid -> CH0_TIME_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src22_startofpacket;                                                           // cmd_xbar_demux_001:src22_startofpacket -> CH0_TIME_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] cmd_xbar_demux_001_src22_data;                                                                    // cmd_xbar_demux_001:src22_data -> CH0_TIME_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [98:0] cmd_xbar_demux_001_src22_channel;                                                                 // cmd_xbar_demux_001:src22_channel -> CH0_TIME_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src23_endofpacket;                                                             // cmd_xbar_demux_001:src23_endofpacket -> CH0_YN2_MU_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src23_valid;                                                                   // cmd_xbar_demux_001:src23_valid -> CH0_YN2_MU_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src23_startofpacket;                                                           // cmd_xbar_demux_001:src23_startofpacket -> CH0_YN2_MU_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] cmd_xbar_demux_001_src23_data;                                                                    // cmd_xbar_demux_001:src23_data -> CH0_YN2_MU_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [98:0] cmd_xbar_demux_001_src23_channel;                                                                 // cmd_xbar_demux_001:src23_channel -> CH0_YN2_MU_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src24_endofpacket;                                                             // cmd_xbar_demux_001:src24_endofpacket -> CH0_YN2_ML_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src24_valid;                                                                   // cmd_xbar_demux_001:src24_valid -> CH0_YN2_ML_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src24_startofpacket;                                                           // cmd_xbar_demux_001:src24_startofpacket -> CH0_YN2_ML_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] cmd_xbar_demux_001_src24_data;                                                                    // cmd_xbar_demux_001:src24_data -> CH0_YN2_ML_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [98:0] cmd_xbar_demux_001_src24_channel;                                                                 // cmd_xbar_demux_001:src24_channel -> CH0_YN2_ML_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src25_endofpacket;                                                             // cmd_xbar_demux_001:src25_endofpacket -> CH0_YN2_U_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src25_valid;                                                                   // cmd_xbar_demux_001:src25_valid -> CH0_YN2_U_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src25_startofpacket;                                                           // cmd_xbar_demux_001:src25_startofpacket -> CH0_YN2_U_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] cmd_xbar_demux_001_src25_data;                                                                    // cmd_xbar_demux_001:src25_data -> CH0_YN2_U_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [98:0] cmd_xbar_demux_001_src25_channel;                                                                 // cmd_xbar_demux_001:src25_channel -> CH0_YN2_U_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src26_endofpacket;                                                             // cmd_xbar_demux_001:src26_endofpacket -> CH0_YN2_L_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src26_valid;                                                                   // cmd_xbar_demux_001:src26_valid -> CH0_YN2_L_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src26_startofpacket;                                                           // cmd_xbar_demux_001:src26_startofpacket -> CH0_YN2_L_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] cmd_xbar_demux_001_src26_data;                                                                    // cmd_xbar_demux_001:src26_data -> CH0_YN2_L_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [98:0] cmd_xbar_demux_001_src26_channel;                                                                 // cmd_xbar_demux_001:src26_channel -> CH0_YN2_L_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src27_endofpacket;                                                             // cmd_xbar_demux_001:src27_endofpacket -> CH0_YN3_L_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src27_valid;                                                                   // cmd_xbar_demux_001:src27_valid -> CH0_YN3_L_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src27_startofpacket;                                                           // cmd_xbar_demux_001:src27_startofpacket -> CH0_YN3_L_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] cmd_xbar_demux_001_src27_data;                                                                    // cmd_xbar_demux_001:src27_data -> CH0_YN3_L_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [98:0] cmd_xbar_demux_001_src27_channel;                                                                 // cmd_xbar_demux_001:src27_channel -> CH0_YN3_L_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src28_endofpacket;                                                             // cmd_xbar_demux_001:src28_endofpacket -> CH0_YN3_ML_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src28_valid;                                                                   // cmd_xbar_demux_001:src28_valid -> CH0_YN3_ML_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src28_startofpacket;                                                           // cmd_xbar_demux_001:src28_startofpacket -> CH0_YN3_ML_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] cmd_xbar_demux_001_src28_data;                                                                    // cmd_xbar_demux_001:src28_data -> CH0_YN3_ML_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [98:0] cmd_xbar_demux_001_src28_channel;                                                                 // cmd_xbar_demux_001:src28_channel -> CH0_YN3_ML_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src29_endofpacket;                                                             // cmd_xbar_demux_001:src29_endofpacket -> CH0_YN3_MU_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src29_valid;                                                                   // cmd_xbar_demux_001:src29_valid -> CH0_YN3_MU_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src29_startofpacket;                                                           // cmd_xbar_demux_001:src29_startofpacket -> CH0_YN3_MU_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] cmd_xbar_demux_001_src29_data;                                                                    // cmd_xbar_demux_001:src29_data -> CH0_YN3_MU_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [98:0] cmd_xbar_demux_001_src29_channel;                                                                 // cmd_xbar_demux_001:src29_channel -> CH0_YN3_MU_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src30_endofpacket;                                                             // cmd_xbar_demux_001:src30_endofpacket -> CH0_YN3_U_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src30_valid;                                                                   // cmd_xbar_demux_001:src30_valid -> CH0_YN3_U_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src30_startofpacket;                                                           // cmd_xbar_demux_001:src30_startofpacket -> CH0_YN3_U_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] cmd_xbar_demux_001_src30_data;                                                                    // cmd_xbar_demux_001:src30_data -> CH0_YN3_U_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [98:0] cmd_xbar_demux_001_src30_channel;                                                                 // cmd_xbar_demux_001:src30_channel -> CH0_YN3_U_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src31_endofpacket;                                                             // cmd_xbar_demux_001:src31_endofpacket -> CH1_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src31_valid;                                                                   // cmd_xbar_demux_001:src31_valid -> CH1_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src31_startofpacket;                                                           // cmd_xbar_demux_001:src31_startofpacket -> CH1_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] cmd_xbar_demux_001_src31_data;                                                                    // cmd_xbar_demux_001:src31_data -> CH1_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [98:0] cmd_xbar_demux_001_src31_channel;                                                                 // cmd_xbar_demux_001:src31_channel -> CH1_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src32_endofpacket;                                                             // cmd_xbar_demux_001:src32_endofpacket -> CH1_THRESH_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src32_valid;                                                                   // cmd_xbar_demux_001:src32_valid -> CH1_THRESH_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src32_startofpacket;                                                           // cmd_xbar_demux_001:src32_startofpacket -> CH1_THRESH_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] cmd_xbar_demux_001_src32_data;                                                                    // cmd_xbar_demux_001:src32_data -> CH1_THRESH_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [98:0] cmd_xbar_demux_001_src32_channel;                                                                 // cmd_xbar_demux_001:src32_channel -> CH1_THRESH_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src33_endofpacket;                                                             // cmd_xbar_demux_001:src33_endofpacket -> CH1_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src33_valid;                                                                   // cmd_xbar_demux_001:src33_valid -> CH1_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src33_startofpacket;                                                           // cmd_xbar_demux_001:src33_startofpacket -> CH1_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] cmd_xbar_demux_001_src33_data;                                                                    // cmd_xbar_demux_001:src33_data -> CH1_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [98:0] cmd_xbar_demux_001_src33_channel;                                                                 // cmd_xbar_demux_001:src33_channel -> CH1_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src34_endofpacket;                                                             // cmd_xbar_demux_001:src34_endofpacket -> CH1_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src34_valid;                                                                   // cmd_xbar_demux_001:src34_valid -> CH1_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src34_startofpacket;                                                           // cmd_xbar_demux_001:src34_startofpacket -> CH1_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] cmd_xbar_demux_001_src34_data;                                                                    // cmd_xbar_demux_001:src34_data -> CH1_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [98:0] cmd_xbar_demux_001_src34_channel;                                                                 // cmd_xbar_demux_001:src34_channel -> CH1_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src35_endofpacket;                                                             // cmd_xbar_demux_001:src35_endofpacket -> CH1_TIME_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src35_valid;                                                                   // cmd_xbar_demux_001:src35_valid -> CH1_TIME_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src35_startofpacket;                                                           // cmd_xbar_demux_001:src35_startofpacket -> CH1_TIME_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] cmd_xbar_demux_001_src35_data;                                                                    // cmd_xbar_demux_001:src35_data -> CH1_TIME_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [98:0] cmd_xbar_demux_001_src35_channel;                                                                 // cmd_xbar_demux_001:src35_channel -> CH1_TIME_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src36_endofpacket;                                                             // cmd_xbar_demux_001:src36_endofpacket -> CH1_YN1_U_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src36_valid;                                                                   // cmd_xbar_demux_001:src36_valid -> CH1_YN1_U_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src36_startofpacket;                                                           // cmd_xbar_demux_001:src36_startofpacket -> CH1_YN1_U_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] cmd_xbar_demux_001_src36_data;                                                                    // cmd_xbar_demux_001:src36_data -> CH1_YN1_U_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [98:0] cmd_xbar_demux_001_src36_channel;                                                                 // cmd_xbar_demux_001:src36_channel -> CH1_YN1_U_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src37_endofpacket;                                                             // cmd_xbar_demux_001:src37_endofpacket -> CH1_YN1_MU_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src37_valid;                                                                   // cmd_xbar_demux_001:src37_valid -> CH1_YN1_MU_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src37_startofpacket;                                                           // cmd_xbar_demux_001:src37_startofpacket -> CH1_YN1_MU_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] cmd_xbar_demux_001_src37_data;                                                                    // cmd_xbar_demux_001:src37_data -> CH1_YN1_MU_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [98:0] cmd_xbar_demux_001_src37_channel;                                                                 // cmd_xbar_demux_001:src37_channel -> CH1_YN1_MU_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src38_endofpacket;                                                             // cmd_xbar_demux_001:src38_endofpacket -> CH1_YN1_ML_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src38_valid;                                                                   // cmd_xbar_demux_001:src38_valid -> CH1_YN1_ML_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src38_startofpacket;                                                           // cmd_xbar_demux_001:src38_startofpacket -> CH1_YN1_ML_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] cmd_xbar_demux_001_src38_data;                                                                    // cmd_xbar_demux_001:src38_data -> CH1_YN1_ML_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [98:0] cmd_xbar_demux_001_src38_channel;                                                                 // cmd_xbar_demux_001:src38_channel -> CH1_YN1_ML_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src39_endofpacket;                                                             // cmd_xbar_demux_001:src39_endofpacket -> CH1_YN1_L_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src39_valid;                                                                   // cmd_xbar_demux_001:src39_valid -> CH1_YN1_L_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src39_startofpacket;                                                           // cmd_xbar_demux_001:src39_startofpacket -> CH1_YN1_L_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] cmd_xbar_demux_001_src39_data;                                                                    // cmd_xbar_demux_001:src39_data -> CH1_YN1_L_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [98:0] cmd_xbar_demux_001_src39_channel;                                                                 // cmd_xbar_demux_001:src39_channel -> CH1_YN1_L_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src40_endofpacket;                                                             // cmd_xbar_demux_001:src40_endofpacket -> CH1_YN2_U_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src40_valid;                                                                   // cmd_xbar_demux_001:src40_valid -> CH1_YN2_U_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src40_startofpacket;                                                           // cmd_xbar_demux_001:src40_startofpacket -> CH1_YN2_U_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] cmd_xbar_demux_001_src40_data;                                                                    // cmd_xbar_demux_001:src40_data -> CH1_YN2_U_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [98:0] cmd_xbar_demux_001_src40_channel;                                                                 // cmd_xbar_demux_001:src40_channel -> CH1_YN2_U_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src41_endofpacket;                                                             // cmd_xbar_demux_001:src41_endofpacket -> CH1_YN2_MU_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src41_valid;                                                                   // cmd_xbar_demux_001:src41_valid -> CH1_YN2_MU_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src41_startofpacket;                                                           // cmd_xbar_demux_001:src41_startofpacket -> CH1_YN2_MU_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] cmd_xbar_demux_001_src41_data;                                                                    // cmd_xbar_demux_001:src41_data -> CH1_YN2_MU_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [98:0] cmd_xbar_demux_001_src41_channel;                                                                 // cmd_xbar_demux_001:src41_channel -> CH1_YN2_MU_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src42_endofpacket;                                                             // cmd_xbar_demux_001:src42_endofpacket -> CH1_YN2_ML_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src42_valid;                                                                   // cmd_xbar_demux_001:src42_valid -> CH1_YN2_ML_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src42_startofpacket;                                                           // cmd_xbar_demux_001:src42_startofpacket -> CH1_YN2_ML_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] cmd_xbar_demux_001_src42_data;                                                                    // cmd_xbar_demux_001:src42_data -> CH1_YN2_ML_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [98:0] cmd_xbar_demux_001_src42_channel;                                                                 // cmd_xbar_demux_001:src42_channel -> CH1_YN2_ML_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src43_endofpacket;                                                             // cmd_xbar_demux_001:src43_endofpacket -> CH1_YN2_L_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src43_valid;                                                                   // cmd_xbar_demux_001:src43_valid -> CH1_YN2_L_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src43_startofpacket;                                                           // cmd_xbar_demux_001:src43_startofpacket -> CH1_YN2_L_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] cmd_xbar_demux_001_src43_data;                                                                    // cmd_xbar_demux_001:src43_data -> CH1_YN2_L_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [98:0] cmd_xbar_demux_001_src43_channel;                                                                 // cmd_xbar_demux_001:src43_channel -> CH1_YN2_L_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src44_endofpacket;                                                             // cmd_xbar_demux_001:src44_endofpacket -> CH1_YN3_U_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src44_valid;                                                                   // cmd_xbar_demux_001:src44_valid -> CH1_YN3_U_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src44_startofpacket;                                                           // cmd_xbar_demux_001:src44_startofpacket -> CH1_YN3_U_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] cmd_xbar_demux_001_src44_data;                                                                    // cmd_xbar_demux_001:src44_data -> CH1_YN3_U_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [98:0] cmd_xbar_demux_001_src44_channel;                                                                 // cmd_xbar_demux_001:src44_channel -> CH1_YN3_U_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src45_endofpacket;                                                             // cmd_xbar_demux_001:src45_endofpacket -> CH1_YN3_MU_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src45_valid;                                                                   // cmd_xbar_demux_001:src45_valid -> CH1_YN3_MU_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src45_startofpacket;                                                           // cmd_xbar_demux_001:src45_startofpacket -> CH1_YN3_MU_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] cmd_xbar_demux_001_src45_data;                                                                    // cmd_xbar_demux_001:src45_data -> CH1_YN3_MU_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [98:0] cmd_xbar_demux_001_src45_channel;                                                                 // cmd_xbar_demux_001:src45_channel -> CH1_YN3_MU_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src46_endofpacket;                                                             // cmd_xbar_demux_001:src46_endofpacket -> CH1_YN3_ML_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src46_valid;                                                                   // cmd_xbar_demux_001:src46_valid -> CH1_YN3_ML_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src46_startofpacket;                                                           // cmd_xbar_demux_001:src46_startofpacket -> CH1_YN3_ML_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] cmd_xbar_demux_001_src46_data;                                                                    // cmd_xbar_demux_001:src46_data -> CH1_YN3_ML_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [98:0] cmd_xbar_demux_001_src46_channel;                                                                 // cmd_xbar_demux_001:src46_channel -> CH1_YN3_ML_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src47_endofpacket;                                                             // cmd_xbar_demux_001:src47_endofpacket -> CH1_YN3_L_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src47_valid;                                                                   // cmd_xbar_demux_001:src47_valid -> CH1_YN3_L_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src47_startofpacket;                                                           // cmd_xbar_demux_001:src47_startofpacket -> CH1_YN3_L_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] cmd_xbar_demux_001_src47_data;                                                                    // cmd_xbar_demux_001:src47_data -> CH1_YN3_L_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [98:0] cmd_xbar_demux_001_src47_channel;                                                                 // cmd_xbar_demux_001:src47_channel -> CH1_YN3_L_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src48_endofpacket;                                                             // cmd_xbar_demux_001:src48_endofpacket -> CH2_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src48_valid;                                                                   // cmd_xbar_demux_001:src48_valid -> CH2_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src48_startofpacket;                                                           // cmd_xbar_demux_001:src48_startofpacket -> CH2_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] cmd_xbar_demux_001_src48_data;                                                                    // cmd_xbar_demux_001:src48_data -> CH2_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [98:0] cmd_xbar_demux_001_src48_channel;                                                                 // cmd_xbar_demux_001:src48_channel -> CH2_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src49_endofpacket;                                                             // cmd_xbar_demux_001:src49_endofpacket -> CH2_THRESH_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src49_valid;                                                                   // cmd_xbar_demux_001:src49_valid -> CH2_THRESH_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src49_startofpacket;                                                           // cmd_xbar_demux_001:src49_startofpacket -> CH2_THRESH_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] cmd_xbar_demux_001_src49_data;                                                                    // cmd_xbar_demux_001:src49_data -> CH2_THRESH_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [98:0] cmd_xbar_demux_001_src49_channel;                                                                 // cmd_xbar_demux_001:src49_channel -> CH2_THRESH_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src50_endofpacket;                                                             // cmd_xbar_demux_001:src50_endofpacket -> CH2_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src50_valid;                                                                   // cmd_xbar_demux_001:src50_valid -> CH2_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src50_startofpacket;                                                           // cmd_xbar_demux_001:src50_startofpacket -> CH2_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] cmd_xbar_demux_001_src50_data;                                                                    // cmd_xbar_demux_001:src50_data -> CH2_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [98:0] cmd_xbar_demux_001_src50_channel;                                                                 // cmd_xbar_demux_001:src50_channel -> CH2_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src51_endofpacket;                                                             // cmd_xbar_demux_001:src51_endofpacket -> CH2_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src51_valid;                                                                   // cmd_xbar_demux_001:src51_valid -> CH2_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src51_startofpacket;                                                           // cmd_xbar_demux_001:src51_startofpacket -> CH2_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] cmd_xbar_demux_001_src51_data;                                                                    // cmd_xbar_demux_001:src51_data -> CH2_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [98:0] cmd_xbar_demux_001_src51_channel;                                                                 // cmd_xbar_demux_001:src51_channel -> CH2_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src52_endofpacket;                                                             // cmd_xbar_demux_001:src52_endofpacket -> CH2_TIME_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src52_valid;                                                                   // cmd_xbar_demux_001:src52_valid -> CH2_TIME_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src52_startofpacket;                                                           // cmd_xbar_demux_001:src52_startofpacket -> CH2_TIME_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] cmd_xbar_demux_001_src52_data;                                                                    // cmd_xbar_demux_001:src52_data -> CH2_TIME_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [98:0] cmd_xbar_demux_001_src52_channel;                                                                 // cmd_xbar_demux_001:src52_channel -> CH2_TIME_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src53_endofpacket;                                                             // cmd_xbar_demux_001:src53_endofpacket -> CH2_YN1_U_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src53_valid;                                                                   // cmd_xbar_demux_001:src53_valid -> CH2_YN1_U_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src53_startofpacket;                                                           // cmd_xbar_demux_001:src53_startofpacket -> CH2_YN1_U_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] cmd_xbar_demux_001_src53_data;                                                                    // cmd_xbar_demux_001:src53_data -> CH2_YN1_U_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [98:0] cmd_xbar_demux_001_src53_channel;                                                                 // cmd_xbar_demux_001:src53_channel -> CH2_YN1_U_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src54_endofpacket;                                                             // cmd_xbar_demux_001:src54_endofpacket -> CH2_YN1_MU_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src54_valid;                                                                   // cmd_xbar_demux_001:src54_valid -> CH2_YN1_MU_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src54_startofpacket;                                                           // cmd_xbar_demux_001:src54_startofpacket -> CH2_YN1_MU_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] cmd_xbar_demux_001_src54_data;                                                                    // cmd_xbar_demux_001:src54_data -> CH2_YN1_MU_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [98:0] cmd_xbar_demux_001_src54_channel;                                                                 // cmd_xbar_demux_001:src54_channel -> CH2_YN1_MU_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src55_endofpacket;                                                             // cmd_xbar_demux_001:src55_endofpacket -> CH2_YN1_ML_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src55_valid;                                                                   // cmd_xbar_demux_001:src55_valid -> CH2_YN1_ML_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src55_startofpacket;                                                           // cmd_xbar_demux_001:src55_startofpacket -> CH2_YN1_ML_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] cmd_xbar_demux_001_src55_data;                                                                    // cmd_xbar_demux_001:src55_data -> CH2_YN1_ML_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [98:0] cmd_xbar_demux_001_src55_channel;                                                                 // cmd_xbar_demux_001:src55_channel -> CH2_YN1_ML_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src56_endofpacket;                                                             // cmd_xbar_demux_001:src56_endofpacket -> CH2_YN1_L_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src56_valid;                                                                   // cmd_xbar_demux_001:src56_valid -> CH2_YN1_L_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src56_startofpacket;                                                           // cmd_xbar_demux_001:src56_startofpacket -> CH2_YN1_L_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] cmd_xbar_demux_001_src56_data;                                                                    // cmd_xbar_demux_001:src56_data -> CH2_YN1_L_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [98:0] cmd_xbar_demux_001_src56_channel;                                                                 // cmd_xbar_demux_001:src56_channel -> CH2_YN1_L_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src57_endofpacket;                                                             // cmd_xbar_demux_001:src57_endofpacket -> CH2_YN2_U_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src57_valid;                                                                   // cmd_xbar_demux_001:src57_valid -> CH2_YN2_U_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src57_startofpacket;                                                           // cmd_xbar_demux_001:src57_startofpacket -> CH2_YN2_U_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] cmd_xbar_demux_001_src57_data;                                                                    // cmd_xbar_demux_001:src57_data -> CH2_YN2_U_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [98:0] cmd_xbar_demux_001_src57_channel;                                                                 // cmd_xbar_demux_001:src57_channel -> CH2_YN2_U_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src58_endofpacket;                                                             // cmd_xbar_demux_001:src58_endofpacket -> CH2_YN2_MU_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src58_valid;                                                                   // cmd_xbar_demux_001:src58_valid -> CH2_YN2_MU_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src58_startofpacket;                                                           // cmd_xbar_demux_001:src58_startofpacket -> CH2_YN2_MU_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] cmd_xbar_demux_001_src58_data;                                                                    // cmd_xbar_demux_001:src58_data -> CH2_YN2_MU_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [98:0] cmd_xbar_demux_001_src58_channel;                                                                 // cmd_xbar_demux_001:src58_channel -> CH2_YN2_MU_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src59_endofpacket;                                                             // cmd_xbar_demux_001:src59_endofpacket -> CH2_YN2_ML_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src59_valid;                                                                   // cmd_xbar_demux_001:src59_valid -> CH2_YN2_ML_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src59_startofpacket;                                                           // cmd_xbar_demux_001:src59_startofpacket -> CH2_YN2_ML_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] cmd_xbar_demux_001_src59_data;                                                                    // cmd_xbar_demux_001:src59_data -> CH2_YN2_ML_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [98:0] cmd_xbar_demux_001_src59_channel;                                                                 // cmd_xbar_demux_001:src59_channel -> CH2_YN2_ML_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src60_endofpacket;                                                             // cmd_xbar_demux_001:src60_endofpacket -> CH2_YN2_L_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src60_valid;                                                                   // cmd_xbar_demux_001:src60_valid -> CH2_YN2_L_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src60_startofpacket;                                                           // cmd_xbar_demux_001:src60_startofpacket -> CH2_YN2_L_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] cmd_xbar_demux_001_src60_data;                                                                    // cmd_xbar_demux_001:src60_data -> CH2_YN2_L_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [98:0] cmd_xbar_demux_001_src60_channel;                                                                 // cmd_xbar_demux_001:src60_channel -> CH2_YN2_L_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src61_endofpacket;                                                             // cmd_xbar_demux_001:src61_endofpacket -> CH2_YN3_U_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src61_valid;                                                                   // cmd_xbar_demux_001:src61_valid -> CH2_YN3_U_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src61_startofpacket;                                                           // cmd_xbar_demux_001:src61_startofpacket -> CH2_YN3_U_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] cmd_xbar_demux_001_src61_data;                                                                    // cmd_xbar_demux_001:src61_data -> CH2_YN3_U_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [98:0] cmd_xbar_demux_001_src61_channel;                                                                 // cmd_xbar_demux_001:src61_channel -> CH2_YN3_U_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src62_endofpacket;                                                             // cmd_xbar_demux_001:src62_endofpacket -> CH2_YN3_MU_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src62_valid;                                                                   // cmd_xbar_demux_001:src62_valid -> CH2_YN3_MU_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src62_startofpacket;                                                           // cmd_xbar_demux_001:src62_startofpacket -> CH2_YN3_MU_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] cmd_xbar_demux_001_src62_data;                                                                    // cmd_xbar_demux_001:src62_data -> CH2_YN3_MU_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [98:0] cmd_xbar_demux_001_src62_channel;                                                                 // cmd_xbar_demux_001:src62_channel -> CH2_YN3_MU_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src63_endofpacket;                                                             // cmd_xbar_demux_001:src63_endofpacket -> CH2_YN3_ML_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src63_valid;                                                                   // cmd_xbar_demux_001:src63_valid -> CH2_YN3_ML_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src63_startofpacket;                                                           // cmd_xbar_demux_001:src63_startofpacket -> CH2_YN3_ML_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] cmd_xbar_demux_001_src63_data;                                                                    // cmd_xbar_demux_001:src63_data -> CH2_YN3_ML_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [98:0] cmd_xbar_demux_001_src63_channel;                                                                 // cmd_xbar_demux_001:src63_channel -> CH2_YN3_ML_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src64_endofpacket;                                                             // cmd_xbar_demux_001:src64_endofpacket -> CH2_YN3_L_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src64_valid;                                                                   // cmd_xbar_demux_001:src64_valid -> CH2_YN3_L_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src64_startofpacket;                                                           // cmd_xbar_demux_001:src64_startofpacket -> CH2_YN3_L_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] cmd_xbar_demux_001_src64_data;                                                                    // cmd_xbar_demux_001:src64_data -> CH2_YN3_L_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [98:0] cmd_xbar_demux_001_src64_channel;                                                                 // cmd_xbar_demux_001:src64_channel -> CH2_YN3_L_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src65_endofpacket;                                                             // cmd_xbar_demux_001:src65_endofpacket -> CH3_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src65_valid;                                                                   // cmd_xbar_demux_001:src65_valid -> CH3_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src65_startofpacket;                                                           // cmd_xbar_demux_001:src65_startofpacket -> CH3_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] cmd_xbar_demux_001_src65_data;                                                                    // cmd_xbar_demux_001:src65_data -> CH3_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [98:0] cmd_xbar_demux_001_src65_channel;                                                                 // cmd_xbar_demux_001:src65_channel -> CH3_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src66_endofpacket;                                                             // cmd_xbar_demux_001:src66_endofpacket -> CH3_THRESH_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src66_valid;                                                                   // cmd_xbar_demux_001:src66_valid -> CH3_THRESH_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src66_startofpacket;                                                           // cmd_xbar_demux_001:src66_startofpacket -> CH3_THRESH_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] cmd_xbar_demux_001_src66_data;                                                                    // cmd_xbar_demux_001:src66_data -> CH3_THRESH_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [98:0] cmd_xbar_demux_001_src66_channel;                                                                 // cmd_xbar_demux_001:src66_channel -> CH3_THRESH_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src67_endofpacket;                                                             // cmd_xbar_demux_001:src67_endofpacket -> CH3_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src67_valid;                                                                   // cmd_xbar_demux_001:src67_valid -> CH3_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src67_startofpacket;                                                           // cmd_xbar_demux_001:src67_startofpacket -> CH3_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] cmd_xbar_demux_001_src67_data;                                                                    // cmd_xbar_demux_001:src67_data -> CH3_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [98:0] cmd_xbar_demux_001_src67_channel;                                                                 // cmd_xbar_demux_001:src67_channel -> CH3_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src68_endofpacket;                                                             // cmd_xbar_demux_001:src68_endofpacket -> CH3_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src68_valid;                                                                   // cmd_xbar_demux_001:src68_valid -> CH3_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src68_startofpacket;                                                           // cmd_xbar_demux_001:src68_startofpacket -> CH3_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] cmd_xbar_demux_001_src68_data;                                                                    // cmd_xbar_demux_001:src68_data -> CH3_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [98:0] cmd_xbar_demux_001_src68_channel;                                                                 // cmd_xbar_demux_001:src68_channel -> CH3_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src69_endofpacket;                                                             // cmd_xbar_demux_001:src69_endofpacket -> CH3_YN1_U_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src69_valid;                                                                   // cmd_xbar_demux_001:src69_valid -> CH3_YN1_U_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src69_startofpacket;                                                           // cmd_xbar_demux_001:src69_startofpacket -> CH3_YN1_U_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] cmd_xbar_demux_001_src69_data;                                                                    // cmd_xbar_demux_001:src69_data -> CH3_YN1_U_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [98:0] cmd_xbar_demux_001_src69_channel;                                                                 // cmd_xbar_demux_001:src69_channel -> CH3_YN1_U_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src70_endofpacket;                                                             // cmd_xbar_demux_001:src70_endofpacket -> CH3_TIME_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src70_valid;                                                                   // cmd_xbar_demux_001:src70_valid -> CH3_TIME_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src70_startofpacket;                                                           // cmd_xbar_demux_001:src70_startofpacket -> CH3_TIME_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] cmd_xbar_demux_001_src70_data;                                                                    // cmd_xbar_demux_001:src70_data -> CH3_TIME_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [98:0] cmd_xbar_demux_001_src70_channel;                                                                 // cmd_xbar_demux_001:src70_channel -> CH3_TIME_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src71_endofpacket;                                                             // cmd_xbar_demux_001:src71_endofpacket -> CH3_YN3_L_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src71_valid;                                                                   // cmd_xbar_demux_001:src71_valid -> CH3_YN3_L_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src71_startofpacket;                                                           // cmd_xbar_demux_001:src71_startofpacket -> CH3_YN3_L_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] cmd_xbar_demux_001_src71_data;                                                                    // cmd_xbar_demux_001:src71_data -> CH3_YN3_L_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [98:0] cmd_xbar_demux_001_src71_channel;                                                                 // cmd_xbar_demux_001:src71_channel -> CH3_YN3_L_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src72_endofpacket;                                                             // cmd_xbar_demux_001:src72_endofpacket -> CH3_YN3_ML_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src72_valid;                                                                   // cmd_xbar_demux_001:src72_valid -> CH3_YN3_ML_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src72_startofpacket;                                                           // cmd_xbar_demux_001:src72_startofpacket -> CH3_YN3_ML_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] cmd_xbar_demux_001_src72_data;                                                                    // cmd_xbar_demux_001:src72_data -> CH3_YN3_ML_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [98:0] cmd_xbar_demux_001_src72_channel;                                                                 // cmd_xbar_demux_001:src72_channel -> CH3_YN3_ML_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src73_endofpacket;                                                             // cmd_xbar_demux_001:src73_endofpacket -> CH3_YN3_MU_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src73_valid;                                                                   // cmd_xbar_demux_001:src73_valid -> CH3_YN3_MU_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src73_startofpacket;                                                           // cmd_xbar_demux_001:src73_startofpacket -> CH3_YN3_MU_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] cmd_xbar_demux_001_src73_data;                                                                    // cmd_xbar_demux_001:src73_data -> CH3_YN3_MU_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [98:0] cmd_xbar_demux_001_src73_channel;                                                                 // cmd_xbar_demux_001:src73_channel -> CH3_YN3_MU_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src74_endofpacket;                                                             // cmd_xbar_demux_001:src74_endofpacket -> CH3_YN3_U_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src74_valid;                                                                   // cmd_xbar_demux_001:src74_valid -> CH3_YN3_U_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src74_startofpacket;                                                           // cmd_xbar_demux_001:src74_startofpacket -> CH3_YN3_U_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] cmd_xbar_demux_001_src74_data;                                                                    // cmd_xbar_demux_001:src74_data -> CH3_YN3_U_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [98:0] cmd_xbar_demux_001_src74_channel;                                                                 // cmd_xbar_demux_001:src74_channel -> CH3_YN3_U_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src75_endofpacket;                                                             // cmd_xbar_demux_001:src75_endofpacket -> CH3_YN2_L_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src75_valid;                                                                   // cmd_xbar_demux_001:src75_valid -> CH3_YN2_L_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src75_startofpacket;                                                           // cmd_xbar_demux_001:src75_startofpacket -> CH3_YN2_L_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] cmd_xbar_demux_001_src75_data;                                                                    // cmd_xbar_demux_001:src75_data -> CH3_YN2_L_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [98:0] cmd_xbar_demux_001_src75_channel;                                                                 // cmd_xbar_demux_001:src75_channel -> CH3_YN2_L_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src76_endofpacket;                                                             // cmd_xbar_demux_001:src76_endofpacket -> CH3_YN2_ML_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src76_valid;                                                                   // cmd_xbar_demux_001:src76_valid -> CH3_YN2_ML_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src76_startofpacket;                                                           // cmd_xbar_demux_001:src76_startofpacket -> CH3_YN2_ML_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] cmd_xbar_demux_001_src76_data;                                                                    // cmd_xbar_demux_001:src76_data -> CH3_YN2_ML_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [98:0] cmd_xbar_demux_001_src76_channel;                                                                 // cmd_xbar_demux_001:src76_channel -> CH3_YN2_ML_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src77_endofpacket;                                                             // cmd_xbar_demux_001:src77_endofpacket -> CH3_YN2_MU_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src77_valid;                                                                   // cmd_xbar_demux_001:src77_valid -> CH3_YN2_MU_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src77_startofpacket;                                                           // cmd_xbar_demux_001:src77_startofpacket -> CH3_YN2_MU_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] cmd_xbar_demux_001_src77_data;                                                                    // cmd_xbar_demux_001:src77_data -> CH3_YN2_MU_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [98:0] cmd_xbar_demux_001_src77_channel;                                                                 // cmd_xbar_demux_001:src77_channel -> CH3_YN2_MU_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src78_endofpacket;                                                             // cmd_xbar_demux_001:src78_endofpacket -> CH3_YN2_U_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src78_valid;                                                                   // cmd_xbar_demux_001:src78_valid -> CH3_YN2_U_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src78_startofpacket;                                                           // cmd_xbar_demux_001:src78_startofpacket -> CH3_YN2_U_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] cmd_xbar_demux_001_src78_data;                                                                    // cmd_xbar_demux_001:src78_data -> CH3_YN2_U_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [98:0] cmd_xbar_demux_001_src78_channel;                                                                 // cmd_xbar_demux_001:src78_channel -> CH3_YN2_U_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src79_endofpacket;                                                             // cmd_xbar_demux_001:src79_endofpacket -> CH3_YN1_L_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src79_valid;                                                                   // cmd_xbar_demux_001:src79_valid -> CH3_YN1_L_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src79_startofpacket;                                                           // cmd_xbar_demux_001:src79_startofpacket -> CH3_YN1_L_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] cmd_xbar_demux_001_src79_data;                                                                    // cmd_xbar_demux_001:src79_data -> CH3_YN1_L_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [98:0] cmd_xbar_demux_001_src79_channel;                                                                 // cmd_xbar_demux_001:src79_channel -> CH3_YN1_L_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src80_endofpacket;                                                             // cmd_xbar_demux_001:src80_endofpacket -> CH3_YN1_MU_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src80_valid;                                                                   // cmd_xbar_demux_001:src80_valid -> CH3_YN1_MU_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src80_startofpacket;                                                           // cmd_xbar_demux_001:src80_startofpacket -> CH3_YN1_MU_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] cmd_xbar_demux_001_src80_data;                                                                    // cmd_xbar_demux_001:src80_data -> CH3_YN1_MU_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [98:0] cmd_xbar_demux_001_src80_channel;                                                                 // cmd_xbar_demux_001:src80_channel -> CH3_YN1_MU_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src81_endofpacket;                                                             // cmd_xbar_demux_001:src81_endofpacket -> CH3_YN1_ML_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src81_valid;                                                                   // cmd_xbar_demux_001:src81_valid -> CH3_YN1_ML_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src81_startofpacket;                                                           // cmd_xbar_demux_001:src81_startofpacket -> CH3_YN1_ML_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] cmd_xbar_demux_001_src81_data;                                                                    // cmd_xbar_demux_001:src81_data -> CH3_YN1_ML_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [98:0] cmd_xbar_demux_001_src81_channel;                                                                 // cmd_xbar_demux_001:src81_channel -> CH3_YN1_ML_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src82_endofpacket;                                                             // cmd_xbar_demux_001:src82_endofpacket -> CH4_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src82_valid;                                                                   // cmd_xbar_demux_001:src82_valid -> CH4_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src82_startofpacket;                                                           // cmd_xbar_demux_001:src82_startofpacket -> CH4_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] cmd_xbar_demux_001_src82_data;                                                                    // cmd_xbar_demux_001:src82_data -> CH4_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [98:0] cmd_xbar_demux_001_src82_channel;                                                                 // cmd_xbar_demux_001:src82_channel -> CH4_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src83_endofpacket;                                                             // cmd_xbar_demux_001:src83_endofpacket -> CH4_THRESH_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src83_valid;                                                                   // cmd_xbar_demux_001:src83_valid -> CH4_THRESH_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src83_startofpacket;                                                           // cmd_xbar_demux_001:src83_startofpacket -> CH4_THRESH_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] cmd_xbar_demux_001_src83_data;                                                                    // cmd_xbar_demux_001:src83_data -> CH4_THRESH_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [98:0] cmd_xbar_demux_001_src83_channel;                                                                 // cmd_xbar_demux_001:src83_channel -> CH4_THRESH_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src84_endofpacket;                                                             // cmd_xbar_demux_001:src84_endofpacket -> CH4_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src84_valid;                                                                   // cmd_xbar_demux_001:src84_valid -> CH4_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src84_startofpacket;                                                           // cmd_xbar_demux_001:src84_startofpacket -> CH4_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] cmd_xbar_demux_001_src84_data;                                                                    // cmd_xbar_demux_001:src84_data -> CH4_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [98:0] cmd_xbar_demux_001_src84_channel;                                                                 // cmd_xbar_demux_001:src84_channel -> CH4_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src85_endofpacket;                                                             // cmd_xbar_demux_001:src85_endofpacket -> CH4_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src85_valid;                                                                   // cmd_xbar_demux_001:src85_valid -> CH4_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src85_startofpacket;                                                           // cmd_xbar_demux_001:src85_startofpacket -> CH4_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] cmd_xbar_demux_001_src85_data;                                                                    // cmd_xbar_demux_001:src85_data -> CH4_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [98:0] cmd_xbar_demux_001_src85_channel;                                                                 // cmd_xbar_demux_001:src85_channel -> CH4_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src86_endofpacket;                                                             // cmd_xbar_demux_001:src86_endofpacket -> CH4_TIME_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src86_valid;                                                                   // cmd_xbar_demux_001:src86_valid -> CH4_TIME_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src86_startofpacket;                                                           // cmd_xbar_demux_001:src86_startofpacket -> CH4_TIME_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] cmd_xbar_demux_001_src86_data;                                                                    // cmd_xbar_demux_001:src86_data -> CH4_TIME_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [98:0] cmd_xbar_demux_001_src86_channel;                                                                 // cmd_xbar_demux_001:src86_channel -> CH4_TIME_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src87_endofpacket;                                                             // cmd_xbar_demux_001:src87_endofpacket -> CH4_YN1_U_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src87_valid;                                                                   // cmd_xbar_demux_001:src87_valid -> CH4_YN1_U_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src87_startofpacket;                                                           // cmd_xbar_demux_001:src87_startofpacket -> CH4_YN1_U_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] cmd_xbar_demux_001_src87_data;                                                                    // cmd_xbar_demux_001:src87_data -> CH4_YN1_U_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [98:0] cmd_xbar_demux_001_src87_channel;                                                                 // cmd_xbar_demux_001:src87_channel -> CH4_YN1_U_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src88_endofpacket;                                                             // cmd_xbar_demux_001:src88_endofpacket -> CH4_YN1_MU_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src88_valid;                                                                   // cmd_xbar_demux_001:src88_valid -> CH4_YN1_MU_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src88_startofpacket;                                                           // cmd_xbar_demux_001:src88_startofpacket -> CH4_YN1_MU_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] cmd_xbar_demux_001_src88_data;                                                                    // cmd_xbar_demux_001:src88_data -> CH4_YN1_MU_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [98:0] cmd_xbar_demux_001_src88_channel;                                                                 // cmd_xbar_demux_001:src88_channel -> CH4_YN1_MU_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src89_endofpacket;                                                             // cmd_xbar_demux_001:src89_endofpacket -> CH4_YN1_ML_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src89_valid;                                                                   // cmd_xbar_demux_001:src89_valid -> CH4_YN1_ML_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src89_startofpacket;                                                           // cmd_xbar_demux_001:src89_startofpacket -> CH4_YN1_ML_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] cmd_xbar_demux_001_src89_data;                                                                    // cmd_xbar_demux_001:src89_data -> CH4_YN1_ML_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [98:0] cmd_xbar_demux_001_src89_channel;                                                                 // cmd_xbar_demux_001:src89_channel -> CH4_YN1_ML_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src90_endofpacket;                                                             // cmd_xbar_demux_001:src90_endofpacket -> CH4_YN1_L_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src90_valid;                                                                   // cmd_xbar_demux_001:src90_valid -> CH4_YN1_L_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src90_startofpacket;                                                           // cmd_xbar_demux_001:src90_startofpacket -> CH4_YN1_L_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] cmd_xbar_demux_001_src90_data;                                                                    // cmd_xbar_demux_001:src90_data -> CH4_YN1_L_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [98:0] cmd_xbar_demux_001_src90_channel;                                                                 // cmd_xbar_demux_001:src90_channel -> CH4_YN1_L_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src91_endofpacket;                                                             // cmd_xbar_demux_001:src91_endofpacket -> CH4_YN2_U_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src91_valid;                                                                   // cmd_xbar_demux_001:src91_valid -> CH4_YN2_U_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src91_startofpacket;                                                           // cmd_xbar_demux_001:src91_startofpacket -> CH4_YN2_U_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] cmd_xbar_demux_001_src91_data;                                                                    // cmd_xbar_demux_001:src91_data -> CH4_YN2_U_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [98:0] cmd_xbar_demux_001_src91_channel;                                                                 // cmd_xbar_demux_001:src91_channel -> CH4_YN2_U_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src92_endofpacket;                                                             // cmd_xbar_demux_001:src92_endofpacket -> CH4_YN2_MU_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src92_valid;                                                                   // cmd_xbar_demux_001:src92_valid -> CH4_YN2_MU_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src92_startofpacket;                                                           // cmd_xbar_demux_001:src92_startofpacket -> CH4_YN2_MU_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] cmd_xbar_demux_001_src92_data;                                                                    // cmd_xbar_demux_001:src92_data -> CH4_YN2_MU_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [98:0] cmd_xbar_demux_001_src92_channel;                                                                 // cmd_xbar_demux_001:src92_channel -> CH4_YN2_MU_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src93_endofpacket;                                                             // cmd_xbar_demux_001:src93_endofpacket -> CH4_YN2_ML_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src93_valid;                                                                   // cmd_xbar_demux_001:src93_valid -> CH4_YN2_ML_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src93_startofpacket;                                                           // cmd_xbar_demux_001:src93_startofpacket -> CH4_YN2_ML_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] cmd_xbar_demux_001_src93_data;                                                                    // cmd_xbar_demux_001:src93_data -> CH4_YN2_ML_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [98:0] cmd_xbar_demux_001_src93_channel;                                                                 // cmd_xbar_demux_001:src93_channel -> CH4_YN2_ML_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src94_endofpacket;                                                             // cmd_xbar_demux_001:src94_endofpacket -> CH4_YN2_L_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src94_valid;                                                                   // cmd_xbar_demux_001:src94_valid -> CH4_YN2_L_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src94_startofpacket;                                                           // cmd_xbar_demux_001:src94_startofpacket -> CH4_YN2_L_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] cmd_xbar_demux_001_src94_data;                                                                    // cmd_xbar_demux_001:src94_data -> CH4_YN2_L_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [98:0] cmd_xbar_demux_001_src94_channel;                                                                 // cmd_xbar_demux_001:src94_channel -> CH4_YN2_L_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src95_endofpacket;                                                             // cmd_xbar_demux_001:src95_endofpacket -> CH4_YN3_U_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src95_valid;                                                                   // cmd_xbar_demux_001:src95_valid -> CH4_YN3_U_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src95_startofpacket;                                                           // cmd_xbar_demux_001:src95_startofpacket -> CH4_YN3_U_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] cmd_xbar_demux_001_src95_data;                                                                    // cmd_xbar_demux_001:src95_data -> CH4_YN3_U_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [98:0] cmd_xbar_demux_001_src95_channel;                                                                 // cmd_xbar_demux_001:src95_channel -> CH4_YN3_U_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src96_endofpacket;                                                             // cmd_xbar_demux_001:src96_endofpacket -> CH4_YN3_MU_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src96_valid;                                                                   // cmd_xbar_demux_001:src96_valid -> CH4_YN3_MU_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src96_startofpacket;                                                           // cmd_xbar_demux_001:src96_startofpacket -> CH4_YN3_MU_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] cmd_xbar_demux_001_src96_data;                                                                    // cmd_xbar_demux_001:src96_data -> CH4_YN3_MU_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [98:0] cmd_xbar_demux_001_src96_channel;                                                                 // cmd_xbar_demux_001:src96_channel -> CH4_YN3_MU_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src97_endofpacket;                                                             // cmd_xbar_demux_001:src97_endofpacket -> CH4_YN3_ML_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src97_valid;                                                                   // cmd_xbar_demux_001:src97_valid -> CH4_YN3_ML_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src97_startofpacket;                                                           // cmd_xbar_demux_001:src97_startofpacket -> CH4_YN3_ML_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] cmd_xbar_demux_001_src97_data;                                                                    // cmd_xbar_demux_001:src97_data -> CH4_YN3_ML_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [98:0] cmd_xbar_demux_001_src97_channel;                                                                 // cmd_xbar_demux_001:src97_channel -> CH4_YN3_ML_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src98_endofpacket;                                                             // cmd_xbar_demux_001:src98_endofpacket -> CH4_YN3_L_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src98_valid;                                                                   // cmd_xbar_demux_001:src98_valid -> CH4_YN3_L_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src98_startofpacket;                                                           // cmd_xbar_demux_001:src98_startofpacket -> CH4_YN3_L_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] cmd_xbar_demux_001_src98_data;                                                                    // cmd_xbar_demux_001:src98_data -> CH4_YN3_L_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [98:0] cmd_xbar_demux_001_src98_channel;                                                                 // cmd_xbar_demux_001:src98_channel -> CH4_YN3_L_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          rsp_xbar_demux_src0_endofpacket;                                                                  // rsp_xbar_demux:src0_endofpacket -> rsp_xbar_mux:sink0_endofpacket
	wire          rsp_xbar_demux_src0_valid;                                                                        // rsp_xbar_demux:src0_valid -> rsp_xbar_mux:sink0_valid
	wire          rsp_xbar_demux_src0_startofpacket;                                                                // rsp_xbar_demux:src0_startofpacket -> rsp_xbar_mux:sink0_startofpacket
	wire  [102:0] rsp_xbar_demux_src0_data;                                                                         // rsp_xbar_demux:src0_data -> rsp_xbar_mux:sink0_data
	wire   [98:0] rsp_xbar_demux_src0_channel;                                                                      // rsp_xbar_demux:src0_channel -> rsp_xbar_mux:sink0_channel
	wire          rsp_xbar_demux_src0_ready;                                                                        // rsp_xbar_mux:sink0_ready -> rsp_xbar_demux:src0_ready
	wire          rsp_xbar_demux_src1_endofpacket;                                                                  // rsp_xbar_demux:src1_endofpacket -> rsp_xbar_mux_001:sink0_endofpacket
	wire          rsp_xbar_demux_src1_valid;                                                                        // rsp_xbar_demux:src1_valid -> rsp_xbar_mux_001:sink0_valid
	wire          rsp_xbar_demux_src1_startofpacket;                                                                // rsp_xbar_demux:src1_startofpacket -> rsp_xbar_mux_001:sink0_startofpacket
	wire  [102:0] rsp_xbar_demux_src1_data;                                                                         // rsp_xbar_demux:src1_data -> rsp_xbar_mux_001:sink0_data
	wire   [98:0] rsp_xbar_demux_src1_channel;                                                                      // rsp_xbar_demux:src1_channel -> rsp_xbar_mux_001:sink0_channel
	wire          rsp_xbar_demux_src1_ready;                                                                        // rsp_xbar_mux_001:sink0_ready -> rsp_xbar_demux:src1_ready
	wire          rsp_xbar_demux_001_src0_endofpacket;                                                              // rsp_xbar_demux_001:src0_endofpacket -> rsp_xbar_mux:sink1_endofpacket
	wire          rsp_xbar_demux_001_src0_valid;                                                                    // rsp_xbar_demux_001:src0_valid -> rsp_xbar_mux:sink1_valid
	wire          rsp_xbar_demux_001_src0_startofpacket;                                                            // rsp_xbar_demux_001:src0_startofpacket -> rsp_xbar_mux:sink1_startofpacket
	wire  [102:0] rsp_xbar_demux_001_src0_data;                                                                     // rsp_xbar_demux_001:src0_data -> rsp_xbar_mux:sink1_data
	wire   [98:0] rsp_xbar_demux_001_src0_channel;                                                                  // rsp_xbar_demux_001:src0_channel -> rsp_xbar_mux:sink1_channel
	wire          rsp_xbar_demux_001_src0_ready;                                                                    // rsp_xbar_mux:sink1_ready -> rsp_xbar_demux_001:src0_ready
	wire          rsp_xbar_demux_001_src1_endofpacket;                                                              // rsp_xbar_demux_001:src1_endofpacket -> rsp_xbar_mux_001:sink1_endofpacket
	wire          rsp_xbar_demux_001_src1_valid;                                                                    // rsp_xbar_demux_001:src1_valid -> rsp_xbar_mux_001:sink1_valid
	wire          rsp_xbar_demux_001_src1_startofpacket;                                                            // rsp_xbar_demux_001:src1_startofpacket -> rsp_xbar_mux_001:sink1_startofpacket
	wire  [102:0] rsp_xbar_demux_001_src1_data;                                                                     // rsp_xbar_demux_001:src1_data -> rsp_xbar_mux_001:sink1_data
	wire   [98:0] rsp_xbar_demux_001_src1_channel;                                                                  // rsp_xbar_demux_001:src1_channel -> rsp_xbar_mux_001:sink1_channel
	wire          rsp_xbar_demux_001_src1_ready;                                                                    // rsp_xbar_mux_001:sink1_ready -> rsp_xbar_demux_001:src1_ready
	wire          rsp_xbar_demux_002_src0_endofpacket;                                                              // rsp_xbar_demux_002:src0_endofpacket -> rsp_xbar_mux:sink2_endofpacket
	wire          rsp_xbar_demux_002_src0_valid;                                                                    // rsp_xbar_demux_002:src0_valid -> rsp_xbar_mux:sink2_valid
	wire          rsp_xbar_demux_002_src0_startofpacket;                                                            // rsp_xbar_demux_002:src0_startofpacket -> rsp_xbar_mux:sink2_startofpacket
	wire  [102:0] rsp_xbar_demux_002_src0_data;                                                                     // rsp_xbar_demux_002:src0_data -> rsp_xbar_mux:sink2_data
	wire   [98:0] rsp_xbar_demux_002_src0_channel;                                                                  // rsp_xbar_demux_002:src0_channel -> rsp_xbar_mux:sink2_channel
	wire          rsp_xbar_demux_002_src0_ready;                                                                    // rsp_xbar_mux:sink2_ready -> rsp_xbar_demux_002:src0_ready
	wire          rsp_xbar_demux_002_src1_endofpacket;                                                              // rsp_xbar_demux_002:src1_endofpacket -> rsp_xbar_mux_001:sink2_endofpacket
	wire          rsp_xbar_demux_002_src1_valid;                                                                    // rsp_xbar_demux_002:src1_valid -> rsp_xbar_mux_001:sink2_valid
	wire          rsp_xbar_demux_002_src1_startofpacket;                                                            // rsp_xbar_demux_002:src1_startofpacket -> rsp_xbar_mux_001:sink2_startofpacket
	wire  [102:0] rsp_xbar_demux_002_src1_data;                                                                     // rsp_xbar_demux_002:src1_data -> rsp_xbar_mux_001:sink2_data
	wire   [98:0] rsp_xbar_demux_002_src1_channel;                                                                  // rsp_xbar_demux_002:src1_channel -> rsp_xbar_mux_001:sink2_channel
	wire          rsp_xbar_demux_002_src1_ready;                                                                    // rsp_xbar_mux_001:sink2_ready -> rsp_xbar_demux_002:src1_ready
	wire          rsp_xbar_demux_003_src0_endofpacket;                                                              // rsp_xbar_demux_003:src0_endofpacket -> rsp_xbar_mux_001:sink3_endofpacket
	wire          rsp_xbar_demux_003_src0_valid;                                                                    // rsp_xbar_demux_003:src0_valid -> rsp_xbar_mux_001:sink3_valid
	wire          rsp_xbar_demux_003_src0_startofpacket;                                                            // rsp_xbar_demux_003:src0_startofpacket -> rsp_xbar_mux_001:sink3_startofpacket
	wire  [102:0] rsp_xbar_demux_003_src0_data;                                                                     // rsp_xbar_demux_003:src0_data -> rsp_xbar_mux_001:sink3_data
	wire   [98:0] rsp_xbar_demux_003_src0_channel;                                                                  // rsp_xbar_demux_003:src0_channel -> rsp_xbar_mux_001:sink3_channel
	wire          rsp_xbar_demux_003_src0_ready;                                                                    // rsp_xbar_mux_001:sink3_ready -> rsp_xbar_demux_003:src0_ready
	wire          rsp_xbar_demux_004_src0_endofpacket;                                                              // rsp_xbar_demux_004:src0_endofpacket -> rsp_xbar_mux_001:sink4_endofpacket
	wire          rsp_xbar_demux_004_src0_valid;                                                                    // rsp_xbar_demux_004:src0_valid -> rsp_xbar_mux_001:sink4_valid
	wire          rsp_xbar_demux_004_src0_startofpacket;                                                            // rsp_xbar_demux_004:src0_startofpacket -> rsp_xbar_mux_001:sink4_startofpacket
	wire  [102:0] rsp_xbar_demux_004_src0_data;                                                                     // rsp_xbar_demux_004:src0_data -> rsp_xbar_mux_001:sink4_data
	wire   [98:0] rsp_xbar_demux_004_src0_channel;                                                                  // rsp_xbar_demux_004:src0_channel -> rsp_xbar_mux_001:sink4_channel
	wire          rsp_xbar_demux_004_src0_ready;                                                                    // rsp_xbar_mux_001:sink4_ready -> rsp_xbar_demux_004:src0_ready
	wire          rsp_xbar_demux_005_src0_endofpacket;                                                              // rsp_xbar_demux_005:src0_endofpacket -> rsp_xbar_mux_001:sink5_endofpacket
	wire          rsp_xbar_demux_005_src0_valid;                                                                    // rsp_xbar_demux_005:src0_valid -> rsp_xbar_mux_001:sink5_valid
	wire          rsp_xbar_demux_005_src0_startofpacket;                                                            // rsp_xbar_demux_005:src0_startofpacket -> rsp_xbar_mux_001:sink5_startofpacket
	wire  [102:0] rsp_xbar_demux_005_src0_data;                                                                     // rsp_xbar_demux_005:src0_data -> rsp_xbar_mux_001:sink5_data
	wire   [98:0] rsp_xbar_demux_005_src0_channel;                                                                  // rsp_xbar_demux_005:src0_channel -> rsp_xbar_mux_001:sink5_channel
	wire          rsp_xbar_demux_005_src0_ready;                                                                    // rsp_xbar_mux_001:sink5_ready -> rsp_xbar_demux_005:src0_ready
	wire          rsp_xbar_demux_006_src0_endofpacket;                                                              // rsp_xbar_demux_006:src0_endofpacket -> rsp_xbar_mux_001:sink6_endofpacket
	wire          rsp_xbar_demux_006_src0_valid;                                                                    // rsp_xbar_demux_006:src0_valid -> rsp_xbar_mux_001:sink6_valid
	wire          rsp_xbar_demux_006_src0_startofpacket;                                                            // rsp_xbar_demux_006:src0_startofpacket -> rsp_xbar_mux_001:sink6_startofpacket
	wire  [102:0] rsp_xbar_demux_006_src0_data;                                                                     // rsp_xbar_demux_006:src0_data -> rsp_xbar_mux_001:sink6_data
	wire   [98:0] rsp_xbar_demux_006_src0_channel;                                                                  // rsp_xbar_demux_006:src0_channel -> rsp_xbar_mux_001:sink6_channel
	wire          rsp_xbar_demux_006_src0_ready;                                                                    // rsp_xbar_mux_001:sink6_ready -> rsp_xbar_demux_006:src0_ready
	wire          rsp_xbar_demux_007_src0_endofpacket;                                                              // rsp_xbar_demux_007:src0_endofpacket -> rsp_xbar_mux_001:sink7_endofpacket
	wire          rsp_xbar_demux_007_src0_valid;                                                                    // rsp_xbar_demux_007:src0_valid -> rsp_xbar_mux_001:sink7_valid
	wire          rsp_xbar_demux_007_src0_startofpacket;                                                            // rsp_xbar_demux_007:src0_startofpacket -> rsp_xbar_mux_001:sink7_startofpacket
	wire  [102:0] rsp_xbar_demux_007_src0_data;                                                                     // rsp_xbar_demux_007:src0_data -> rsp_xbar_mux_001:sink7_data
	wire   [98:0] rsp_xbar_demux_007_src0_channel;                                                                  // rsp_xbar_demux_007:src0_channel -> rsp_xbar_mux_001:sink7_channel
	wire          rsp_xbar_demux_007_src0_ready;                                                                    // rsp_xbar_mux_001:sink7_ready -> rsp_xbar_demux_007:src0_ready
	wire          rsp_xbar_demux_008_src0_endofpacket;                                                              // rsp_xbar_demux_008:src0_endofpacket -> rsp_xbar_mux_001:sink8_endofpacket
	wire          rsp_xbar_demux_008_src0_valid;                                                                    // rsp_xbar_demux_008:src0_valid -> rsp_xbar_mux_001:sink8_valid
	wire          rsp_xbar_demux_008_src0_startofpacket;                                                            // rsp_xbar_demux_008:src0_startofpacket -> rsp_xbar_mux_001:sink8_startofpacket
	wire  [102:0] rsp_xbar_demux_008_src0_data;                                                                     // rsp_xbar_demux_008:src0_data -> rsp_xbar_mux_001:sink8_data
	wire   [98:0] rsp_xbar_demux_008_src0_channel;                                                                  // rsp_xbar_demux_008:src0_channel -> rsp_xbar_mux_001:sink8_channel
	wire          rsp_xbar_demux_008_src0_ready;                                                                    // rsp_xbar_mux_001:sink8_ready -> rsp_xbar_demux_008:src0_ready
	wire          rsp_xbar_demux_009_src0_endofpacket;                                                              // rsp_xbar_demux_009:src0_endofpacket -> rsp_xbar_mux_001:sink9_endofpacket
	wire          rsp_xbar_demux_009_src0_valid;                                                                    // rsp_xbar_demux_009:src0_valid -> rsp_xbar_mux_001:sink9_valid
	wire          rsp_xbar_demux_009_src0_startofpacket;                                                            // rsp_xbar_demux_009:src0_startofpacket -> rsp_xbar_mux_001:sink9_startofpacket
	wire  [102:0] rsp_xbar_demux_009_src0_data;                                                                     // rsp_xbar_demux_009:src0_data -> rsp_xbar_mux_001:sink9_data
	wire   [98:0] rsp_xbar_demux_009_src0_channel;                                                                  // rsp_xbar_demux_009:src0_channel -> rsp_xbar_mux_001:sink9_channel
	wire          rsp_xbar_demux_009_src0_ready;                                                                    // rsp_xbar_mux_001:sink9_ready -> rsp_xbar_demux_009:src0_ready
	wire          rsp_xbar_demux_010_src0_endofpacket;                                                              // rsp_xbar_demux_010:src0_endofpacket -> rsp_xbar_mux_001:sink10_endofpacket
	wire          rsp_xbar_demux_010_src0_valid;                                                                    // rsp_xbar_demux_010:src0_valid -> rsp_xbar_mux_001:sink10_valid
	wire          rsp_xbar_demux_010_src0_startofpacket;                                                            // rsp_xbar_demux_010:src0_startofpacket -> rsp_xbar_mux_001:sink10_startofpacket
	wire  [102:0] rsp_xbar_demux_010_src0_data;                                                                     // rsp_xbar_demux_010:src0_data -> rsp_xbar_mux_001:sink10_data
	wire   [98:0] rsp_xbar_demux_010_src0_channel;                                                                  // rsp_xbar_demux_010:src0_channel -> rsp_xbar_mux_001:sink10_channel
	wire          rsp_xbar_demux_010_src0_ready;                                                                    // rsp_xbar_mux_001:sink10_ready -> rsp_xbar_demux_010:src0_ready
	wire          rsp_xbar_demux_011_src0_endofpacket;                                                              // rsp_xbar_demux_011:src0_endofpacket -> rsp_xbar_mux_001:sink11_endofpacket
	wire          rsp_xbar_demux_011_src0_valid;                                                                    // rsp_xbar_demux_011:src0_valid -> rsp_xbar_mux_001:sink11_valid
	wire          rsp_xbar_demux_011_src0_startofpacket;                                                            // rsp_xbar_demux_011:src0_startofpacket -> rsp_xbar_mux_001:sink11_startofpacket
	wire  [102:0] rsp_xbar_demux_011_src0_data;                                                                     // rsp_xbar_demux_011:src0_data -> rsp_xbar_mux_001:sink11_data
	wire   [98:0] rsp_xbar_demux_011_src0_channel;                                                                  // rsp_xbar_demux_011:src0_channel -> rsp_xbar_mux_001:sink11_channel
	wire          rsp_xbar_demux_011_src0_ready;                                                                    // rsp_xbar_mux_001:sink11_ready -> rsp_xbar_demux_011:src0_ready
	wire          rsp_xbar_demux_012_src0_endofpacket;                                                              // rsp_xbar_demux_012:src0_endofpacket -> rsp_xbar_mux_001:sink12_endofpacket
	wire          rsp_xbar_demux_012_src0_valid;                                                                    // rsp_xbar_demux_012:src0_valid -> rsp_xbar_mux_001:sink12_valid
	wire          rsp_xbar_demux_012_src0_startofpacket;                                                            // rsp_xbar_demux_012:src0_startofpacket -> rsp_xbar_mux_001:sink12_startofpacket
	wire  [102:0] rsp_xbar_demux_012_src0_data;                                                                     // rsp_xbar_demux_012:src0_data -> rsp_xbar_mux_001:sink12_data
	wire   [98:0] rsp_xbar_demux_012_src0_channel;                                                                  // rsp_xbar_demux_012:src0_channel -> rsp_xbar_mux_001:sink12_channel
	wire          rsp_xbar_demux_012_src0_ready;                                                                    // rsp_xbar_mux_001:sink12_ready -> rsp_xbar_demux_012:src0_ready
	wire          rsp_xbar_demux_013_src0_endofpacket;                                                              // rsp_xbar_demux_013:src0_endofpacket -> rsp_xbar_mux_001:sink13_endofpacket
	wire          rsp_xbar_demux_013_src0_valid;                                                                    // rsp_xbar_demux_013:src0_valid -> rsp_xbar_mux_001:sink13_valid
	wire          rsp_xbar_demux_013_src0_startofpacket;                                                            // rsp_xbar_demux_013:src0_startofpacket -> rsp_xbar_mux_001:sink13_startofpacket
	wire  [102:0] rsp_xbar_demux_013_src0_data;                                                                     // rsp_xbar_demux_013:src0_data -> rsp_xbar_mux_001:sink13_data
	wire   [98:0] rsp_xbar_demux_013_src0_channel;                                                                  // rsp_xbar_demux_013:src0_channel -> rsp_xbar_mux_001:sink13_channel
	wire          rsp_xbar_demux_013_src0_ready;                                                                    // rsp_xbar_mux_001:sink13_ready -> rsp_xbar_demux_013:src0_ready
	wire          rsp_xbar_demux_014_src0_endofpacket;                                                              // rsp_xbar_demux_014:src0_endofpacket -> rsp_xbar_mux_001:sink14_endofpacket
	wire          rsp_xbar_demux_014_src0_valid;                                                                    // rsp_xbar_demux_014:src0_valid -> rsp_xbar_mux_001:sink14_valid
	wire          rsp_xbar_demux_014_src0_startofpacket;                                                            // rsp_xbar_demux_014:src0_startofpacket -> rsp_xbar_mux_001:sink14_startofpacket
	wire  [102:0] rsp_xbar_demux_014_src0_data;                                                                     // rsp_xbar_demux_014:src0_data -> rsp_xbar_mux_001:sink14_data
	wire   [98:0] rsp_xbar_demux_014_src0_channel;                                                                  // rsp_xbar_demux_014:src0_channel -> rsp_xbar_mux_001:sink14_channel
	wire          rsp_xbar_demux_014_src0_ready;                                                                    // rsp_xbar_mux_001:sink14_ready -> rsp_xbar_demux_014:src0_ready
	wire          rsp_xbar_demux_015_src0_endofpacket;                                                              // rsp_xbar_demux_015:src0_endofpacket -> rsp_xbar_mux_001:sink15_endofpacket
	wire          rsp_xbar_demux_015_src0_valid;                                                                    // rsp_xbar_demux_015:src0_valid -> rsp_xbar_mux_001:sink15_valid
	wire          rsp_xbar_demux_015_src0_startofpacket;                                                            // rsp_xbar_demux_015:src0_startofpacket -> rsp_xbar_mux_001:sink15_startofpacket
	wire  [102:0] rsp_xbar_demux_015_src0_data;                                                                     // rsp_xbar_demux_015:src0_data -> rsp_xbar_mux_001:sink15_data
	wire   [98:0] rsp_xbar_demux_015_src0_channel;                                                                  // rsp_xbar_demux_015:src0_channel -> rsp_xbar_mux_001:sink15_channel
	wire          rsp_xbar_demux_015_src0_ready;                                                                    // rsp_xbar_mux_001:sink15_ready -> rsp_xbar_demux_015:src0_ready
	wire          rsp_xbar_demux_016_src0_endofpacket;                                                              // rsp_xbar_demux_016:src0_endofpacket -> rsp_xbar_mux_001:sink16_endofpacket
	wire          rsp_xbar_demux_016_src0_valid;                                                                    // rsp_xbar_demux_016:src0_valid -> rsp_xbar_mux_001:sink16_valid
	wire          rsp_xbar_demux_016_src0_startofpacket;                                                            // rsp_xbar_demux_016:src0_startofpacket -> rsp_xbar_mux_001:sink16_startofpacket
	wire  [102:0] rsp_xbar_demux_016_src0_data;                                                                     // rsp_xbar_demux_016:src0_data -> rsp_xbar_mux_001:sink16_data
	wire   [98:0] rsp_xbar_demux_016_src0_channel;                                                                  // rsp_xbar_demux_016:src0_channel -> rsp_xbar_mux_001:sink16_channel
	wire          rsp_xbar_demux_016_src0_ready;                                                                    // rsp_xbar_mux_001:sink16_ready -> rsp_xbar_demux_016:src0_ready
	wire          rsp_xbar_demux_017_src0_endofpacket;                                                              // rsp_xbar_demux_017:src0_endofpacket -> rsp_xbar_mux_001:sink17_endofpacket
	wire          rsp_xbar_demux_017_src0_valid;                                                                    // rsp_xbar_demux_017:src0_valid -> rsp_xbar_mux_001:sink17_valid
	wire          rsp_xbar_demux_017_src0_startofpacket;                                                            // rsp_xbar_demux_017:src0_startofpacket -> rsp_xbar_mux_001:sink17_startofpacket
	wire  [102:0] rsp_xbar_demux_017_src0_data;                                                                     // rsp_xbar_demux_017:src0_data -> rsp_xbar_mux_001:sink17_data
	wire   [98:0] rsp_xbar_demux_017_src0_channel;                                                                  // rsp_xbar_demux_017:src0_channel -> rsp_xbar_mux_001:sink17_channel
	wire          rsp_xbar_demux_017_src0_ready;                                                                    // rsp_xbar_mux_001:sink17_ready -> rsp_xbar_demux_017:src0_ready
	wire          rsp_xbar_demux_018_src0_endofpacket;                                                              // rsp_xbar_demux_018:src0_endofpacket -> rsp_xbar_mux_001:sink18_endofpacket
	wire          rsp_xbar_demux_018_src0_valid;                                                                    // rsp_xbar_demux_018:src0_valid -> rsp_xbar_mux_001:sink18_valid
	wire          rsp_xbar_demux_018_src0_startofpacket;                                                            // rsp_xbar_demux_018:src0_startofpacket -> rsp_xbar_mux_001:sink18_startofpacket
	wire  [102:0] rsp_xbar_demux_018_src0_data;                                                                     // rsp_xbar_demux_018:src0_data -> rsp_xbar_mux_001:sink18_data
	wire   [98:0] rsp_xbar_demux_018_src0_channel;                                                                  // rsp_xbar_demux_018:src0_channel -> rsp_xbar_mux_001:sink18_channel
	wire          rsp_xbar_demux_018_src0_ready;                                                                    // rsp_xbar_mux_001:sink18_ready -> rsp_xbar_demux_018:src0_ready
	wire          rsp_xbar_demux_019_src0_endofpacket;                                                              // rsp_xbar_demux_019:src0_endofpacket -> rsp_xbar_mux_001:sink19_endofpacket
	wire          rsp_xbar_demux_019_src0_valid;                                                                    // rsp_xbar_demux_019:src0_valid -> rsp_xbar_mux_001:sink19_valid
	wire          rsp_xbar_demux_019_src0_startofpacket;                                                            // rsp_xbar_demux_019:src0_startofpacket -> rsp_xbar_mux_001:sink19_startofpacket
	wire  [102:0] rsp_xbar_demux_019_src0_data;                                                                     // rsp_xbar_demux_019:src0_data -> rsp_xbar_mux_001:sink19_data
	wire   [98:0] rsp_xbar_demux_019_src0_channel;                                                                  // rsp_xbar_demux_019:src0_channel -> rsp_xbar_mux_001:sink19_channel
	wire          rsp_xbar_demux_019_src0_ready;                                                                    // rsp_xbar_mux_001:sink19_ready -> rsp_xbar_demux_019:src0_ready
	wire          rsp_xbar_demux_020_src0_endofpacket;                                                              // rsp_xbar_demux_020:src0_endofpacket -> rsp_xbar_mux_001:sink20_endofpacket
	wire          rsp_xbar_demux_020_src0_valid;                                                                    // rsp_xbar_demux_020:src0_valid -> rsp_xbar_mux_001:sink20_valid
	wire          rsp_xbar_demux_020_src0_startofpacket;                                                            // rsp_xbar_demux_020:src0_startofpacket -> rsp_xbar_mux_001:sink20_startofpacket
	wire  [102:0] rsp_xbar_demux_020_src0_data;                                                                     // rsp_xbar_demux_020:src0_data -> rsp_xbar_mux_001:sink20_data
	wire   [98:0] rsp_xbar_demux_020_src0_channel;                                                                  // rsp_xbar_demux_020:src0_channel -> rsp_xbar_mux_001:sink20_channel
	wire          rsp_xbar_demux_020_src0_ready;                                                                    // rsp_xbar_mux_001:sink20_ready -> rsp_xbar_demux_020:src0_ready
	wire          rsp_xbar_demux_021_src0_endofpacket;                                                              // rsp_xbar_demux_021:src0_endofpacket -> rsp_xbar_mux_001:sink21_endofpacket
	wire          rsp_xbar_demux_021_src0_valid;                                                                    // rsp_xbar_demux_021:src0_valid -> rsp_xbar_mux_001:sink21_valid
	wire          rsp_xbar_demux_021_src0_startofpacket;                                                            // rsp_xbar_demux_021:src0_startofpacket -> rsp_xbar_mux_001:sink21_startofpacket
	wire  [102:0] rsp_xbar_demux_021_src0_data;                                                                     // rsp_xbar_demux_021:src0_data -> rsp_xbar_mux_001:sink21_data
	wire   [98:0] rsp_xbar_demux_021_src0_channel;                                                                  // rsp_xbar_demux_021:src0_channel -> rsp_xbar_mux_001:sink21_channel
	wire          rsp_xbar_demux_021_src0_ready;                                                                    // rsp_xbar_mux_001:sink21_ready -> rsp_xbar_demux_021:src0_ready
	wire          rsp_xbar_demux_022_src0_endofpacket;                                                              // rsp_xbar_demux_022:src0_endofpacket -> rsp_xbar_mux_001:sink22_endofpacket
	wire          rsp_xbar_demux_022_src0_valid;                                                                    // rsp_xbar_demux_022:src0_valid -> rsp_xbar_mux_001:sink22_valid
	wire          rsp_xbar_demux_022_src0_startofpacket;                                                            // rsp_xbar_demux_022:src0_startofpacket -> rsp_xbar_mux_001:sink22_startofpacket
	wire  [102:0] rsp_xbar_demux_022_src0_data;                                                                     // rsp_xbar_demux_022:src0_data -> rsp_xbar_mux_001:sink22_data
	wire   [98:0] rsp_xbar_demux_022_src0_channel;                                                                  // rsp_xbar_demux_022:src0_channel -> rsp_xbar_mux_001:sink22_channel
	wire          rsp_xbar_demux_022_src0_ready;                                                                    // rsp_xbar_mux_001:sink22_ready -> rsp_xbar_demux_022:src0_ready
	wire          rsp_xbar_demux_023_src0_endofpacket;                                                              // rsp_xbar_demux_023:src0_endofpacket -> rsp_xbar_mux_001:sink23_endofpacket
	wire          rsp_xbar_demux_023_src0_valid;                                                                    // rsp_xbar_demux_023:src0_valid -> rsp_xbar_mux_001:sink23_valid
	wire          rsp_xbar_demux_023_src0_startofpacket;                                                            // rsp_xbar_demux_023:src0_startofpacket -> rsp_xbar_mux_001:sink23_startofpacket
	wire  [102:0] rsp_xbar_demux_023_src0_data;                                                                     // rsp_xbar_demux_023:src0_data -> rsp_xbar_mux_001:sink23_data
	wire   [98:0] rsp_xbar_demux_023_src0_channel;                                                                  // rsp_xbar_demux_023:src0_channel -> rsp_xbar_mux_001:sink23_channel
	wire          rsp_xbar_demux_023_src0_ready;                                                                    // rsp_xbar_mux_001:sink23_ready -> rsp_xbar_demux_023:src0_ready
	wire          rsp_xbar_demux_024_src0_endofpacket;                                                              // rsp_xbar_demux_024:src0_endofpacket -> rsp_xbar_mux_001:sink24_endofpacket
	wire          rsp_xbar_demux_024_src0_valid;                                                                    // rsp_xbar_demux_024:src0_valid -> rsp_xbar_mux_001:sink24_valid
	wire          rsp_xbar_demux_024_src0_startofpacket;                                                            // rsp_xbar_demux_024:src0_startofpacket -> rsp_xbar_mux_001:sink24_startofpacket
	wire  [102:0] rsp_xbar_demux_024_src0_data;                                                                     // rsp_xbar_demux_024:src0_data -> rsp_xbar_mux_001:sink24_data
	wire   [98:0] rsp_xbar_demux_024_src0_channel;                                                                  // rsp_xbar_demux_024:src0_channel -> rsp_xbar_mux_001:sink24_channel
	wire          rsp_xbar_demux_024_src0_ready;                                                                    // rsp_xbar_mux_001:sink24_ready -> rsp_xbar_demux_024:src0_ready
	wire          rsp_xbar_demux_025_src0_endofpacket;                                                              // rsp_xbar_demux_025:src0_endofpacket -> rsp_xbar_mux_001:sink25_endofpacket
	wire          rsp_xbar_demux_025_src0_valid;                                                                    // rsp_xbar_demux_025:src0_valid -> rsp_xbar_mux_001:sink25_valid
	wire          rsp_xbar_demux_025_src0_startofpacket;                                                            // rsp_xbar_demux_025:src0_startofpacket -> rsp_xbar_mux_001:sink25_startofpacket
	wire  [102:0] rsp_xbar_demux_025_src0_data;                                                                     // rsp_xbar_demux_025:src0_data -> rsp_xbar_mux_001:sink25_data
	wire   [98:0] rsp_xbar_demux_025_src0_channel;                                                                  // rsp_xbar_demux_025:src0_channel -> rsp_xbar_mux_001:sink25_channel
	wire          rsp_xbar_demux_025_src0_ready;                                                                    // rsp_xbar_mux_001:sink25_ready -> rsp_xbar_demux_025:src0_ready
	wire          rsp_xbar_demux_026_src0_endofpacket;                                                              // rsp_xbar_demux_026:src0_endofpacket -> rsp_xbar_mux_001:sink26_endofpacket
	wire          rsp_xbar_demux_026_src0_valid;                                                                    // rsp_xbar_demux_026:src0_valid -> rsp_xbar_mux_001:sink26_valid
	wire          rsp_xbar_demux_026_src0_startofpacket;                                                            // rsp_xbar_demux_026:src0_startofpacket -> rsp_xbar_mux_001:sink26_startofpacket
	wire  [102:0] rsp_xbar_demux_026_src0_data;                                                                     // rsp_xbar_demux_026:src0_data -> rsp_xbar_mux_001:sink26_data
	wire   [98:0] rsp_xbar_demux_026_src0_channel;                                                                  // rsp_xbar_demux_026:src0_channel -> rsp_xbar_mux_001:sink26_channel
	wire          rsp_xbar_demux_026_src0_ready;                                                                    // rsp_xbar_mux_001:sink26_ready -> rsp_xbar_demux_026:src0_ready
	wire          rsp_xbar_demux_027_src0_endofpacket;                                                              // rsp_xbar_demux_027:src0_endofpacket -> rsp_xbar_mux_001:sink27_endofpacket
	wire          rsp_xbar_demux_027_src0_valid;                                                                    // rsp_xbar_demux_027:src0_valid -> rsp_xbar_mux_001:sink27_valid
	wire          rsp_xbar_demux_027_src0_startofpacket;                                                            // rsp_xbar_demux_027:src0_startofpacket -> rsp_xbar_mux_001:sink27_startofpacket
	wire  [102:0] rsp_xbar_demux_027_src0_data;                                                                     // rsp_xbar_demux_027:src0_data -> rsp_xbar_mux_001:sink27_data
	wire   [98:0] rsp_xbar_demux_027_src0_channel;                                                                  // rsp_xbar_demux_027:src0_channel -> rsp_xbar_mux_001:sink27_channel
	wire          rsp_xbar_demux_027_src0_ready;                                                                    // rsp_xbar_mux_001:sink27_ready -> rsp_xbar_demux_027:src0_ready
	wire          rsp_xbar_demux_028_src0_endofpacket;                                                              // rsp_xbar_demux_028:src0_endofpacket -> rsp_xbar_mux_001:sink28_endofpacket
	wire          rsp_xbar_demux_028_src0_valid;                                                                    // rsp_xbar_demux_028:src0_valid -> rsp_xbar_mux_001:sink28_valid
	wire          rsp_xbar_demux_028_src0_startofpacket;                                                            // rsp_xbar_demux_028:src0_startofpacket -> rsp_xbar_mux_001:sink28_startofpacket
	wire  [102:0] rsp_xbar_demux_028_src0_data;                                                                     // rsp_xbar_demux_028:src0_data -> rsp_xbar_mux_001:sink28_data
	wire   [98:0] rsp_xbar_demux_028_src0_channel;                                                                  // rsp_xbar_demux_028:src0_channel -> rsp_xbar_mux_001:sink28_channel
	wire          rsp_xbar_demux_028_src0_ready;                                                                    // rsp_xbar_mux_001:sink28_ready -> rsp_xbar_demux_028:src0_ready
	wire          rsp_xbar_demux_029_src0_endofpacket;                                                              // rsp_xbar_demux_029:src0_endofpacket -> rsp_xbar_mux_001:sink29_endofpacket
	wire          rsp_xbar_demux_029_src0_valid;                                                                    // rsp_xbar_demux_029:src0_valid -> rsp_xbar_mux_001:sink29_valid
	wire          rsp_xbar_demux_029_src0_startofpacket;                                                            // rsp_xbar_demux_029:src0_startofpacket -> rsp_xbar_mux_001:sink29_startofpacket
	wire  [102:0] rsp_xbar_demux_029_src0_data;                                                                     // rsp_xbar_demux_029:src0_data -> rsp_xbar_mux_001:sink29_data
	wire   [98:0] rsp_xbar_demux_029_src0_channel;                                                                  // rsp_xbar_demux_029:src0_channel -> rsp_xbar_mux_001:sink29_channel
	wire          rsp_xbar_demux_029_src0_ready;                                                                    // rsp_xbar_mux_001:sink29_ready -> rsp_xbar_demux_029:src0_ready
	wire          rsp_xbar_demux_030_src0_endofpacket;                                                              // rsp_xbar_demux_030:src0_endofpacket -> rsp_xbar_mux_001:sink30_endofpacket
	wire          rsp_xbar_demux_030_src0_valid;                                                                    // rsp_xbar_demux_030:src0_valid -> rsp_xbar_mux_001:sink30_valid
	wire          rsp_xbar_demux_030_src0_startofpacket;                                                            // rsp_xbar_demux_030:src0_startofpacket -> rsp_xbar_mux_001:sink30_startofpacket
	wire  [102:0] rsp_xbar_demux_030_src0_data;                                                                     // rsp_xbar_demux_030:src0_data -> rsp_xbar_mux_001:sink30_data
	wire   [98:0] rsp_xbar_demux_030_src0_channel;                                                                  // rsp_xbar_demux_030:src0_channel -> rsp_xbar_mux_001:sink30_channel
	wire          rsp_xbar_demux_030_src0_ready;                                                                    // rsp_xbar_mux_001:sink30_ready -> rsp_xbar_demux_030:src0_ready
	wire          rsp_xbar_demux_031_src0_endofpacket;                                                              // rsp_xbar_demux_031:src0_endofpacket -> rsp_xbar_mux_001:sink31_endofpacket
	wire          rsp_xbar_demux_031_src0_valid;                                                                    // rsp_xbar_demux_031:src0_valid -> rsp_xbar_mux_001:sink31_valid
	wire          rsp_xbar_demux_031_src0_startofpacket;                                                            // rsp_xbar_demux_031:src0_startofpacket -> rsp_xbar_mux_001:sink31_startofpacket
	wire  [102:0] rsp_xbar_demux_031_src0_data;                                                                     // rsp_xbar_demux_031:src0_data -> rsp_xbar_mux_001:sink31_data
	wire   [98:0] rsp_xbar_demux_031_src0_channel;                                                                  // rsp_xbar_demux_031:src0_channel -> rsp_xbar_mux_001:sink31_channel
	wire          rsp_xbar_demux_031_src0_ready;                                                                    // rsp_xbar_mux_001:sink31_ready -> rsp_xbar_demux_031:src0_ready
	wire          rsp_xbar_demux_032_src0_endofpacket;                                                              // rsp_xbar_demux_032:src0_endofpacket -> rsp_xbar_mux_001:sink32_endofpacket
	wire          rsp_xbar_demux_032_src0_valid;                                                                    // rsp_xbar_demux_032:src0_valid -> rsp_xbar_mux_001:sink32_valid
	wire          rsp_xbar_demux_032_src0_startofpacket;                                                            // rsp_xbar_demux_032:src0_startofpacket -> rsp_xbar_mux_001:sink32_startofpacket
	wire  [102:0] rsp_xbar_demux_032_src0_data;                                                                     // rsp_xbar_demux_032:src0_data -> rsp_xbar_mux_001:sink32_data
	wire   [98:0] rsp_xbar_demux_032_src0_channel;                                                                  // rsp_xbar_demux_032:src0_channel -> rsp_xbar_mux_001:sink32_channel
	wire          rsp_xbar_demux_032_src0_ready;                                                                    // rsp_xbar_mux_001:sink32_ready -> rsp_xbar_demux_032:src0_ready
	wire          rsp_xbar_demux_033_src0_endofpacket;                                                              // rsp_xbar_demux_033:src0_endofpacket -> rsp_xbar_mux_001:sink33_endofpacket
	wire          rsp_xbar_demux_033_src0_valid;                                                                    // rsp_xbar_demux_033:src0_valid -> rsp_xbar_mux_001:sink33_valid
	wire          rsp_xbar_demux_033_src0_startofpacket;                                                            // rsp_xbar_demux_033:src0_startofpacket -> rsp_xbar_mux_001:sink33_startofpacket
	wire  [102:0] rsp_xbar_demux_033_src0_data;                                                                     // rsp_xbar_demux_033:src0_data -> rsp_xbar_mux_001:sink33_data
	wire   [98:0] rsp_xbar_demux_033_src0_channel;                                                                  // rsp_xbar_demux_033:src0_channel -> rsp_xbar_mux_001:sink33_channel
	wire          rsp_xbar_demux_033_src0_ready;                                                                    // rsp_xbar_mux_001:sink33_ready -> rsp_xbar_demux_033:src0_ready
	wire          rsp_xbar_demux_034_src0_endofpacket;                                                              // rsp_xbar_demux_034:src0_endofpacket -> rsp_xbar_mux_001:sink34_endofpacket
	wire          rsp_xbar_demux_034_src0_valid;                                                                    // rsp_xbar_demux_034:src0_valid -> rsp_xbar_mux_001:sink34_valid
	wire          rsp_xbar_demux_034_src0_startofpacket;                                                            // rsp_xbar_demux_034:src0_startofpacket -> rsp_xbar_mux_001:sink34_startofpacket
	wire  [102:0] rsp_xbar_demux_034_src0_data;                                                                     // rsp_xbar_demux_034:src0_data -> rsp_xbar_mux_001:sink34_data
	wire   [98:0] rsp_xbar_demux_034_src0_channel;                                                                  // rsp_xbar_demux_034:src0_channel -> rsp_xbar_mux_001:sink34_channel
	wire          rsp_xbar_demux_034_src0_ready;                                                                    // rsp_xbar_mux_001:sink34_ready -> rsp_xbar_demux_034:src0_ready
	wire          rsp_xbar_demux_035_src0_endofpacket;                                                              // rsp_xbar_demux_035:src0_endofpacket -> rsp_xbar_mux_001:sink35_endofpacket
	wire          rsp_xbar_demux_035_src0_valid;                                                                    // rsp_xbar_demux_035:src0_valid -> rsp_xbar_mux_001:sink35_valid
	wire          rsp_xbar_demux_035_src0_startofpacket;                                                            // rsp_xbar_demux_035:src0_startofpacket -> rsp_xbar_mux_001:sink35_startofpacket
	wire  [102:0] rsp_xbar_demux_035_src0_data;                                                                     // rsp_xbar_demux_035:src0_data -> rsp_xbar_mux_001:sink35_data
	wire   [98:0] rsp_xbar_demux_035_src0_channel;                                                                  // rsp_xbar_demux_035:src0_channel -> rsp_xbar_mux_001:sink35_channel
	wire          rsp_xbar_demux_035_src0_ready;                                                                    // rsp_xbar_mux_001:sink35_ready -> rsp_xbar_demux_035:src0_ready
	wire          rsp_xbar_demux_036_src0_endofpacket;                                                              // rsp_xbar_demux_036:src0_endofpacket -> rsp_xbar_mux_001:sink36_endofpacket
	wire          rsp_xbar_demux_036_src0_valid;                                                                    // rsp_xbar_demux_036:src0_valid -> rsp_xbar_mux_001:sink36_valid
	wire          rsp_xbar_demux_036_src0_startofpacket;                                                            // rsp_xbar_demux_036:src0_startofpacket -> rsp_xbar_mux_001:sink36_startofpacket
	wire  [102:0] rsp_xbar_demux_036_src0_data;                                                                     // rsp_xbar_demux_036:src0_data -> rsp_xbar_mux_001:sink36_data
	wire   [98:0] rsp_xbar_demux_036_src0_channel;                                                                  // rsp_xbar_demux_036:src0_channel -> rsp_xbar_mux_001:sink36_channel
	wire          rsp_xbar_demux_036_src0_ready;                                                                    // rsp_xbar_mux_001:sink36_ready -> rsp_xbar_demux_036:src0_ready
	wire          rsp_xbar_demux_037_src0_endofpacket;                                                              // rsp_xbar_demux_037:src0_endofpacket -> rsp_xbar_mux_001:sink37_endofpacket
	wire          rsp_xbar_demux_037_src0_valid;                                                                    // rsp_xbar_demux_037:src0_valid -> rsp_xbar_mux_001:sink37_valid
	wire          rsp_xbar_demux_037_src0_startofpacket;                                                            // rsp_xbar_demux_037:src0_startofpacket -> rsp_xbar_mux_001:sink37_startofpacket
	wire  [102:0] rsp_xbar_demux_037_src0_data;                                                                     // rsp_xbar_demux_037:src0_data -> rsp_xbar_mux_001:sink37_data
	wire   [98:0] rsp_xbar_demux_037_src0_channel;                                                                  // rsp_xbar_demux_037:src0_channel -> rsp_xbar_mux_001:sink37_channel
	wire          rsp_xbar_demux_037_src0_ready;                                                                    // rsp_xbar_mux_001:sink37_ready -> rsp_xbar_demux_037:src0_ready
	wire          rsp_xbar_demux_038_src0_endofpacket;                                                              // rsp_xbar_demux_038:src0_endofpacket -> rsp_xbar_mux_001:sink38_endofpacket
	wire          rsp_xbar_demux_038_src0_valid;                                                                    // rsp_xbar_demux_038:src0_valid -> rsp_xbar_mux_001:sink38_valid
	wire          rsp_xbar_demux_038_src0_startofpacket;                                                            // rsp_xbar_demux_038:src0_startofpacket -> rsp_xbar_mux_001:sink38_startofpacket
	wire  [102:0] rsp_xbar_demux_038_src0_data;                                                                     // rsp_xbar_demux_038:src0_data -> rsp_xbar_mux_001:sink38_data
	wire   [98:0] rsp_xbar_demux_038_src0_channel;                                                                  // rsp_xbar_demux_038:src0_channel -> rsp_xbar_mux_001:sink38_channel
	wire          rsp_xbar_demux_038_src0_ready;                                                                    // rsp_xbar_mux_001:sink38_ready -> rsp_xbar_demux_038:src0_ready
	wire          rsp_xbar_demux_039_src0_endofpacket;                                                              // rsp_xbar_demux_039:src0_endofpacket -> rsp_xbar_mux_001:sink39_endofpacket
	wire          rsp_xbar_demux_039_src0_valid;                                                                    // rsp_xbar_demux_039:src0_valid -> rsp_xbar_mux_001:sink39_valid
	wire          rsp_xbar_demux_039_src0_startofpacket;                                                            // rsp_xbar_demux_039:src0_startofpacket -> rsp_xbar_mux_001:sink39_startofpacket
	wire  [102:0] rsp_xbar_demux_039_src0_data;                                                                     // rsp_xbar_demux_039:src0_data -> rsp_xbar_mux_001:sink39_data
	wire   [98:0] rsp_xbar_demux_039_src0_channel;                                                                  // rsp_xbar_demux_039:src0_channel -> rsp_xbar_mux_001:sink39_channel
	wire          rsp_xbar_demux_039_src0_ready;                                                                    // rsp_xbar_mux_001:sink39_ready -> rsp_xbar_demux_039:src0_ready
	wire          rsp_xbar_demux_040_src0_endofpacket;                                                              // rsp_xbar_demux_040:src0_endofpacket -> rsp_xbar_mux_001:sink40_endofpacket
	wire          rsp_xbar_demux_040_src0_valid;                                                                    // rsp_xbar_demux_040:src0_valid -> rsp_xbar_mux_001:sink40_valid
	wire          rsp_xbar_demux_040_src0_startofpacket;                                                            // rsp_xbar_demux_040:src0_startofpacket -> rsp_xbar_mux_001:sink40_startofpacket
	wire  [102:0] rsp_xbar_demux_040_src0_data;                                                                     // rsp_xbar_demux_040:src0_data -> rsp_xbar_mux_001:sink40_data
	wire   [98:0] rsp_xbar_demux_040_src0_channel;                                                                  // rsp_xbar_demux_040:src0_channel -> rsp_xbar_mux_001:sink40_channel
	wire          rsp_xbar_demux_040_src0_ready;                                                                    // rsp_xbar_mux_001:sink40_ready -> rsp_xbar_demux_040:src0_ready
	wire          rsp_xbar_demux_041_src0_endofpacket;                                                              // rsp_xbar_demux_041:src0_endofpacket -> rsp_xbar_mux_001:sink41_endofpacket
	wire          rsp_xbar_demux_041_src0_valid;                                                                    // rsp_xbar_demux_041:src0_valid -> rsp_xbar_mux_001:sink41_valid
	wire          rsp_xbar_demux_041_src0_startofpacket;                                                            // rsp_xbar_demux_041:src0_startofpacket -> rsp_xbar_mux_001:sink41_startofpacket
	wire  [102:0] rsp_xbar_demux_041_src0_data;                                                                     // rsp_xbar_demux_041:src0_data -> rsp_xbar_mux_001:sink41_data
	wire   [98:0] rsp_xbar_demux_041_src0_channel;                                                                  // rsp_xbar_demux_041:src0_channel -> rsp_xbar_mux_001:sink41_channel
	wire          rsp_xbar_demux_041_src0_ready;                                                                    // rsp_xbar_mux_001:sink41_ready -> rsp_xbar_demux_041:src0_ready
	wire          rsp_xbar_demux_042_src0_endofpacket;                                                              // rsp_xbar_demux_042:src0_endofpacket -> rsp_xbar_mux_001:sink42_endofpacket
	wire          rsp_xbar_demux_042_src0_valid;                                                                    // rsp_xbar_demux_042:src0_valid -> rsp_xbar_mux_001:sink42_valid
	wire          rsp_xbar_demux_042_src0_startofpacket;                                                            // rsp_xbar_demux_042:src0_startofpacket -> rsp_xbar_mux_001:sink42_startofpacket
	wire  [102:0] rsp_xbar_demux_042_src0_data;                                                                     // rsp_xbar_demux_042:src0_data -> rsp_xbar_mux_001:sink42_data
	wire   [98:0] rsp_xbar_demux_042_src0_channel;                                                                  // rsp_xbar_demux_042:src0_channel -> rsp_xbar_mux_001:sink42_channel
	wire          rsp_xbar_demux_042_src0_ready;                                                                    // rsp_xbar_mux_001:sink42_ready -> rsp_xbar_demux_042:src0_ready
	wire          rsp_xbar_demux_043_src0_endofpacket;                                                              // rsp_xbar_demux_043:src0_endofpacket -> rsp_xbar_mux_001:sink43_endofpacket
	wire          rsp_xbar_demux_043_src0_valid;                                                                    // rsp_xbar_demux_043:src0_valid -> rsp_xbar_mux_001:sink43_valid
	wire          rsp_xbar_demux_043_src0_startofpacket;                                                            // rsp_xbar_demux_043:src0_startofpacket -> rsp_xbar_mux_001:sink43_startofpacket
	wire  [102:0] rsp_xbar_demux_043_src0_data;                                                                     // rsp_xbar_demux_043:src0_data -> rsp_xbar_mux_001:sink43_data
	wire   [98:0] rsp_xbar_demux_043_src0_channel;                                                                  // rsp_xbar_demux_043:src0_channel -> rsp_xbar_mux_001:sink43_channel
	wire          rsp_xbar_demux_043_src0_ready;                                                                    // rsp_xbar_mux_001:sink43_ready -> rsp_xbar_demux_043:src0_ready
	wire          rsp_xbar_demux_044_src0_endofpacket;                                                              // rsp_xbar_demux_044:src0_endofpacket -> rsp_xbar_mux_001:sink44_endofpacket
	wire          rsp_xbar_demux_044_src0_valid;                                                                    // rsp_xbar_demux_044:src0_valid -> rsp_xbar_mux_001:sink44_valid
	wire          rsp_xbar_demux_044_src0_startofpacket;                                                            // rsp_xbar_demux_044:src0_startofpacket -> rsp_xbar_mux_001:sink44_startofpacket
	wire  [102:0] rsp_xbar_demux_044_src0_data;                                                                     // rsp_xbar_demux_044:src0_data -> rsp_xbar_mux_001:sink44_data
	wire   [98:0] rsp_xbar_demux_044_src0_channel;                                                                  // rsp_xbar_demux_044:src0_channel -> rsp_xbar_mux_001:sink44_channel
	wire          rsp_xbar_demux_044_src0_ready;                                                                    // rsp_xbar_mux_001:sink44_ready -> rsp_xbar_demux_044:src0_ready
	wire          rsp_xbar_demux_045_src0_endofpacket;                                                              // rsp_xbar_demux_045:src0_endofpacket -> rsp_xbar_mux_001:sink45_endofpacket
	wire          rsp_xbar_demux_045_src0_valid;                                                                    // rsp_xbar_demux_045:src0_valid -> rsp_xbar_mux_001:sink45_valid
	wire          rsp_xbar_demux_045_src0_startofpacket;                                                            // rsp_xbar_demux_045:src0_startofpacket -> rsp_xbar_mux_001:sink45_startofpacket
	wire  [102:0] rsp_xbar_demux_045_src0_data;                                                                     // rsp_xbar_demux_045:src0_data -> rsp_xbar_mux_001:sink45_data
	wire   [98:0] rsp_xbar_demux_045_src0_channel;                                                                  // rsp_xbar_demux_045:src0_channel -> rsp_xbar_mux_001:sink45_channel
	wire          rsp_xbar_demux_045_src0_ready;                                                                    // rsp_xbar_mux_001:sink45_ready -> rsp_xbar_demux_045:src0_ready
	wire          rsp_xbar_demux_046_src0_endofpacket;                                                              // rsp_xbar_demux_046:src0_endofpacket -> rsp_xbar_mux_001:sink46_endofpacket
	wire          rsp_xbar_demux_046_src0_valid;                                                                    // rsp_xbar_demux_046:src0_valid -> rsp_xbar_mux_001:sink46_valid
	wire          rsp_xbar_demux_046_src0_startofpacket;                                                            // rsp_xbar_demux_046:src0_startofpacket -> rsp_xbar_mux_001:sink46_startofpacket
	wire  [102:0] rsp_xbar_demux_046_src0_data;                                                                     // rsp_xbar_demux_046:src0_data -> rsp_xbar_mux_001:sink46_data
	wire   [98:0] rsp_xbar_demux_046_src0_channel;                                                                  // rsp_xbar_demux_046:src0_channel -> rsp_xbar_mux_001:sink46_channel
	wire          rsp_xbar_demux_046_src0_ready;                                                                    // rsp_xbar_mux_001:sink46_ready -> rsp_xbar_demux_046:src0_ready
	wire          rsp_xbar_demux_047_src0_endofpacket;                                                              // rsp_xbar_demux_047:src0_endofpacket -> rsp_xbar_mux_001:sink47_endofpacket
	wire          rsp_xbar_demux_047_src0_valid;                                                                    // rsp_xbar_demux_047:src0_valid -> rsp_xbar_mux_001:sink47_valid
	wire          rsp_xbar_demux_047_src0_startofpacket;                                                            // rsp_xbar_demux_047:src0_startofpacket -> rsp_xbar_mux_001:sink47_startofpacket
	wire  [102:0] rsp_xbar_demux_047_src0_data;                                                                     // rsp_xbar_demux_047:src0_data -> rsp_xbar_mux_001:sink47_data
	wire   [98:0] rsp_xbar_demux_047_src0_channel;                                                                  // rsp_xbar_demux_047:src0_channel -> rsp_xbar_mux_001:sink47_channel
	wire          rsp_xbar_demux_047_src0_ready;                                                                    // rsp_xbar_mux_001:sink47_ready -> rsp_xbar_demux_047:src0_ready
	wire          rsp_xbar_demux_048_src0_endofpacket;                                                              // rsp_xbar_demux_048:src0_endofpacket -> rsp_xbar_mux_001:sink48_endofpacket
	wire          rsp_xbar_demux_048_src0_valid;                                                                    // rsp_xbar_demux_048:src0_valid -> rsp_xbar_mux_001:sink48_valid
	wire          rsp_xbar_demux_048_src0_startofpacket;                                                            // rsp_xbar_demux_048:src0_startofpacket -> rsp_xbar_mux_001:sink48_startofpacket
	wire  [102:0] rsp_xbar_demux_048_src0_data;                                                                     // rsp_xbar_demux_048:src0_data -> rsp_xbar_mux_001:sink48_data
	wire   [98:0] rsp_xbar_demux_048_src0_channel;                                                                  // rsp_xbar_demux_048:src0_channel -> rsp_xbar_mux_001:sink48_channel
	wire          rsp_xbar_demux_048_src0_ready;                                                                    // rsp_xbar_mux_001:sink48_ready -> rsp_xbar_demux_048:src0_ready
	wire          rsp_xbar_demux_049_src0_endofpacket;                                                              // rsp_xbar_demux_049:src0_endofpacket -> rsp_xbar_mux_001:sink49_endofpacket
	wire          rsp_xbar_demux_049_src0_valid;                                                                    // rsp_xbar_demux_049:src0_valid -> rsp_xbar_mux_001:sink49_valid
	wire          rsp_xbar_demux_049_src0_startofpacket;                                                            // rsp_xbar_demux_049:src0_startofpacket -> rsp_xbar_mux_001:sink49_startofpacket
	wire  [102:0] rsp_xbar_demux_049_src0_data;                                                                     // rsp_xbar_demux_049:src0_data -> rsp_xbar_mux_001:sink49_data
	wire   [98:0] rsp_xbar_demux_049_src0_channel;                                                                  // rsp_xbar_demux_049:src0_channel -> rsp_xbar_mux_001:sink49_channel
	wire          rsp_xbar_demux_049_src0_ready;                                                                    // rsp_xbar_mux_001:sink49_ready -> rsp_xbar_demux_049:src0_ready
	wire          rsp_xbar_demux_050_src0_endofpacket;                                                              // rsp_xbar_demux_050:src0_endofpacket -> rsp_xbar_mux_001:sink50_endofpacket
	wire          rsp_xbar_demux_050_src0_valid;                                                                    // rsp_xbar_demux_050:src0_valid -> rsp_xbar_mux_001:sink50_valid
	wire          rsp_xbar_demux_050_src0_startofpacket;                                                            // rsp_xbar_demux_050:src0_startofpacket -> rsp_xbar_mux_001:sink50_startofpacket
	wire  [102:0] rsp_xbar_demux_050_src0_data;                                                                     // rsp_xbar_demux_050:src0_data -> rsp_xbar_mux_001:sink50_data
	wire   [98:0] rsp_xbar_demux_050_src0_channel;                                                                  // rsp_xbar_demux_050:src0_channel -> rsp_xbar_mux_001:sink50_channel
	wire          rsp_xbar_demux_050_src0_ready;                                                                    // rsp_xbar_mux_001:sink50_ready -> rsp_xbar_demux_050:src0_ready
	wire          rsp_xbar_demux_051_src0_endofpacket;                                                              // rsp_xbar_demux_051:src0_endofpacket -> rsp_xbar_mux_001:sink51_endofpacket
	wire          rsp_xbar_demux_051_src0_valid;                                                                    // rsp_xbar_demux_051:src0_valid -> rsp_xbar_mux_001:sink51_valid
	wire          rsp_xbar_demux_051_src0_startofpacket;                                                            // rsp_xbar_demux_051:src0_startofpacket -> rsp_xbar_mux_001:sink51_startofpacket
	wire  [102:0] rsp_xbar_demux_051_src0_data;                                                                     // rsp_xbar_demux_051:src0_data -> rsp_xbar_mux_001:sink51_data
	wire   [98:0] rsp_xbar_demux_051_src0_channel;                                                                  // rsp_xbar_demux_051:src0_channel -> rsp_xbar_mux_001:sink51_channel
	wire          rsp_xbar_demux_051_src0_ready;                                                                    // rsp_xbar_mux_001:sink51_ready -> rsp_xbar_demux_051:src0_ready
	wire          rsp_xbar_demux_052_src0_endofpacket;                                                              // rsp_xbar_demux_052:src0_endofpacket -> rsp_xbar_mux_001:sink52_endofpacket
	wire          rsp_xbar_demux_052_src0_valid;                                                                    // rsp_xbar_demux_052:src0_valid -> rsp_xbar_mux_001:sink52_valid
	wire          rsp_xbar_demux_052_src0_startofpacket;                                                            // rsp_xbar_demux_052:src0_startofpacket -> rsp_xbar_mux_001:sink52_startofpacket
	wire  [102:0] rsp_xbar_demux_052_src0_data;                                                                     // rsp_xbar_demux_052:src0_data -> rsp_xbar_mux_001:sink52_data
	wire   [98:0] rsp_xbar_demux_052_src0_channel;                                                                  // rsp_xbar_demux_052:src0_channel -> rsp_xbar_mux_001:sink52_channel
	wire          rsp_xbar_demux_052_src0_ready;                                                                    // rsp_xbar_mux_001:sink52_ready -> rsp_xbar_demux_052:src0_ready
	wire          rsp_xbar_demux_053_src0_endofpacket;                                                              // rsp_xbar_demux_053:src0_endofpacket -> rsp_xbar_mux_001:sink53_endofpacket
	wire          rsp_xbar_demux_053_src0_valid;                                                                    // rsp_xbar_demux_053:src0_valid -> rsp_xbar_mux_001:sink53_valid
	wire          rsp_xbar_demux_053_src0_startofpacket;                                                            // rsp_xbar_demux_053:src0_startofpacket -> rsp_xbar_mux_001:sink53_startofpacket
	wire  [102:0] rsp_xbar_demux_053_src0_data;                                                                     // rsp_xbar_demux_053:src0_data -> rsp_xbar_mux_001:sink53_data
	wire   [98:0] rsp_xbar_demux_053_src0_channel;                                                                  // rsp_xbar_demux_053:src0_channel -> rsp_xbar_mux_001:sink53_channel
	wire          rsp_xbar_demux_053_src0_ready;                                                                    // rsp_xbar_mux_001:sink53_ready -> rsp_xbar_demux_053:src0_ready
	wire          rsp_xbar_demux_054_src0_endofpacket;                                                              // rsp_xbar_demux_054:src0_endofpacket -> rsp_xbar_mux_001:sink54_endofpacket
	wire          rsp_xbar_demux_054_src0_valid;                                                                    // rsp_xbar_demux_054:src0_valid -> rsp_xbar_mux_001:sink54_valid
	wire          rsp_xbar_demux_054_src0_startofpacket;                                                            // rsp_xbar_demux_054:src0_startofpacket -> rsp_xbar_mux_001:sink54_startofpacket
	wire  [102:0] rsp_xbar_demux_054_src0_data;                                                                     // rsp_xbar_demux_054:src0_data -> rsp_xbar_mux_001:sink54_data
	wire   [98:0] rsp_xbar_demux_054_src0_channel;                                                                  // rsp_xbar_demux_054:src0_channel -> rsp_xbar_mux_001:sink54_channel
	wire          rsp_xbar_demux_054_src0_ready;                                                                    // rsp_xbar_mux_001:sink54_ready -> rsp_xbar_demux_054:src0_ready
	wire          rsp_xbar_demux_055_src0_endofpacket;                                                              // rsp_xbar_demux_055:src0_endofpacket -> rsp_xbar_mux_001:sink55_endofpacket
	wire          rsp_xbar_demux_055_src0_valid;                                                                    // rsp_xbar_demux_055:src0_valid -> rsp_xbar_mux_001:sink55_valid
	wire          rsp_xbar_demux_055_src0_startofpacket;                                                            // rsp_xbar_demux_055:src0_startofpacket -> rsp_xbar_mux_001:sink55_startofpacket
	wire  [102:0] rsp_xbar_demux_055_src0_data;                                                                     // rsp_xbar_demux_055:src0_data -> rsp_xbar_mux_001:sink55_data
	wire   [98:0] rsp_xbar_demux_055_src0_channel;                                                                  // rsp_xbar_demux_055:src0_channel -> rsp_xbar_mux_001:sink55_channel
	wire          rsp_xbar_demux_055_src0_ready;                                                                    // rsp_xbar_mux_001:sink55_ready -> rsp_xbar_demux_055:src0_ready
	wire          rsp_xbar_demux_056_src0_endofpacket;                                                              // rsp_xbar_demux_056:src0_endofpacket -> rsp_xbar_mux_001:sink56_endofpacket
	wire          rsp_xbar_demux_056_src0_valid;                                                                    // rsp_xbar_demux_056:src0_valid -> rsp_xbar_mux_001:sink56_valid
	wire          rsp_xbar_demux_056_src0_startofpacket;                                                            // rsp_xbar_demux_056:src0_startofpacket -> rsp_xbar_mux_001:sink56_startofpacket
	wire  [102:0] rsp_xbar_demux_056_src0_data;                                                                     // rsp_xbar_demux_056:src0_data -> rsp_xbar_mux_001:sink56_data
	wire   [98:0] rsp_xbar_demux_056_src0_channel;                                                                  // rsp_xbar_demux_056:src0_channel -> rsp_xbar_mux_001:sink56_channel
	wire          rsp_xbar_demux_056_src0_ready;                                                                    // rsp_xbar_mux_001:sink56_ready -> rsp_xbar_demux_056:src0_ready
	wire          rsp_xbar_demux_057_src0_endofpacket;                                                              // rsp_xbar_demux_057:src0_endofpacket -> rsp_xbar_mux_001:sink57_endofpacket
	wire          rsp_xbar_demux_057_src0_valid;                                                                    // rsp_xbar_demux_057:src0_valid -> rsp_xbar_mux_001:sink57_valid
	wire          rsp_xbar_demux_057_src0_startofpacket;                                                            // rsp_xbar_demux_057:src0_startofpacket -> rsp_xbar_mux_001:sink57_startofpacket
	wire  [102:0] rsp_xbar_demux_057_src0_data;                                                                     // rsp_xbar_demux_057:src0_data -> rsp_xbar_mux_001:sink57_data
	wire   [98:0] rsp_xbar_demux_057_src0_channel;                                                                  // rsp_xbar_demux_057:src0_channel -> rsp_xbar_mux_001:sink57_channel
	wire          rsp_xbar_demux_057_src0_ready;                                                                    // rsp_xbar_mux_001:sink57_ready -> rsp_xbar_demux_057:src0_ready
	wire          rsp_xbar_demux_058_src0_endofpacket;                                                              // rsp_xbar_demux_058:src0_endofpacket -> rsp_xbar_mux_001:sink58_endofpacket
	wire          rsp_xbar_demux_058_src0_valid;                                                                    // rsp_xbar_demux_058:src0_valid -> rsp_xbar_mux_001:sink58_valid
	wire          rsp_xbar_demux_058_src0_startofpacket;                                                            // rsp_xbar_demux_058:src0_startofpacket -> rsp_xbar_mux_001:sink58_startofpacket
	wire  [102:0] rsp_xbar_demux_058_src0_data;                                                                     // rsp_xbar_demux_058:src0_data -> rsp_xbar_mux_001:sink58_data
	wire   [98:0] rsp_xbar_demux_058_src0_channel;                                                                  // rsp_xbar_demux_058:src0_channel -> rsp_xbar_mux_001:sink58_channel
	wire          rsp_xbar_demux_058_src0_ready;                                                                    // rsp_xbar_mux_001:sink58_ready -> rsp_xbar_demux_058:src0_ready
	wire          rsp_xbar_demux_059_src0_endofpacket;                                                              // rsp_xbar_demux_059:src0_endofpacket -> rsp_xbar_mux_001:sink59_endofpacket
	wire          rsp_xbar_demux_059_src0_valid;                                                                    // rsp_xbar_demux_059:src0_valid -> rsp_xbar_mux_001:sink59_valid
	wire          rsp_xbar_demux_059_src0_startofpacket;                                                            // rsp_xbar_demux_059:src0_startofpacket -> rsp_xbar_mux_001:sink59_startofpacket
	wire  [102:0] rsp_xbar_demux_059_src0_data;                                                                     // rsp_xbar_demux_059:src0_data -> rsp_xbar_mux_001:sink59_data
	wire   [98:0] rsp_xbar_demux_059_src0_channel;                                                                  // rsp_xbar_demux_059:src0_channel -> rsp_xbar_mux_001:sink59_channel
	wire          rsp_xbar_demux_059_src0_ready;                                                                    // rsp_xbar_mux_001:sink59_ready -> rsp_xbar_demux_059:src0_ready
	wire          rsp_xbar_demux_060_src0_endofpacket;                                                              // rsp_xbar_demux_060:src0_endofpacket -> rsp_xbar_mux_001:sink60_endofpacket
	wire          rsp_xbar_demux_060_src0_valid;                                                                    // rsp_xbar_demux_060:src0_valid -> rsp_xbar_mux_001:sink60_valid
	wire          rsp_xbar_demux_060_src0_startofpacket;                                                            // rsp_xbar_demux_060:src0_startofpacket -> rsp_xbar_mux_001:sink60_startofpacket
	wire  [102:0] rsp_xbar_demux_060_src0_data;                                                                     // rsp_xbar_demux_060:src0_data -> rsp_xbar_mux_001:sink60_data
	wire   [98:0] rsp_xbar_demux_060_src0_channel;                                                                  // rsp_xbar_demux_060:src0_channel -> rsp_xbar_mux_001:sink60_channel
	wire          rsp_xbar_demux_060_src0_ready;                                                                    // rsp_xbar_mux_001:sink60_ready -> rsp_xbar_demux_060:src0_ready
	wire          rsp_xbar_demux_061_src0_endofpacket;                                                              // rsp_xbar_demux_061:src0_endofpacket -> rsp_xbar_mux_001:sink61_endofpacket
	wire          rsp_xbar_demux_061_src0_valid;                                                                    // rsp_xbar_demux_061:src0_valid -> rsp_xbar_mux_001:sink61_valid
	wire          rsp_xbar_demux_061_src0_startofpacket;                                                            // rsp_xbar_demux_061:src0_startofpacket -> rsp_xbar_mux_001:sink61_startofpacket
	wire  [102:0] rsp_xbar_demux_061_src0_data;                                                                     // rsp_xbar_demux_061:src0_data -> rsp_xbar_mux_001:sink61_data
	wire   [98:0] rsp_xbar_demux_061_src0_channel;                                                                  // rsp_xbar_demux_061:src0_channel -> rsp_xbar_mux_001:sink61_channel
	wire          rsp_xbar_demux_061_src0_ready;                                                                    // rsp_xbar_mux_001:sink61_ready -> rsp_xbar_demux_061:src0_ready
	wire          rsp_xbar_demux_062_src0_endofpacket;                                                              // rsp_xbar_demux_062:src0_endofpacket -> rsp_xbar_mux_001:sink62_endofpacket
	wire          rsp_xbar_demux_062_src0_valid;                                                                    // rsp_xbar_demux_062:src0_valid -> rsp_xbar_mux_001:sink62_valid
	wire          rsp_xbar_demux_062_src0_startofpacket;                                                            // rsp_xbar_demux_062:src0_startofpacket -> rsp_xbar_mux_001:sink62_startofpacket
	wire  [102:0] rsp_xbar_demux_062_src0_data;                                                                     // rsp_xbar_demux_062:src0_data -> rsp_xbar_mux_001:sink62_data
	wire   [98:0] rsp_xbar_demux_062_src0_channel;                                                                  // rsp_xbar_demux_062:src0_channel -> rsp_xbar_mux_001:sink62_channel
	wire          rsp_xbar_demux_062_src0_ready;                                                                    // rsp_xbar_mux_001:sink62_ready -> rsp_xbar_demux_062:src0_ready
	wire          rsp_xbar_demux_063_src0_endofpacket;                                                              // rsp_xbar_demux_063:src0_endofpacket -> rsp_xbar_mux_001:sink63_endofpacket
	wire          rsp_xbar_demux_063_src0_valid;                                                                    // rsp_xbar_demux_063:src0_valid -> rsp_xbar_mux_001:sink63_valid
	wire          rsp_xbar_demux_063_src0_startofpacket;                                                            // rsp_xbar_demux_063:src0_startofpacket -> rsp_xbar_mux_001:sink63_startofpacket
	wire  [102:0] rsp_xbar_demux_063_src0_data;                                                                     // rsp_xbar_demux_063:src0_data -> rsp_xbar_mux_001:sink63_data
	wire   [98:0] rsp_xbar_demux_063_src0_channel;                                                                  // rsp_xbar_demux_063:src0_channel -> rsp_xbar_mux_001:sink63_channel
	wire          rsp_xbar_demux_063_src0_ready;                                                                    // rsp_xbar_mux_001:sink63_ready -> rsp_xbar_demux_063:src0_ready
	wire          rsp_xbar_demux_064_src0_endofpacket;                                                              // rsp_xbar_demux_064:src0_endofpacket -> rsp_xbar_mux_001:sink64_endofpacket
	wire          rsp_xbar_demux_064_src0_valid;                                                                    // rsp_xbar_demux_064:src0_valid -> rsp_xbar_mux_001:sink64_valid
	wire          rsp_xbar_demux_064_src0_startofpacket;                                                            // rsp_xbar_demux_064:src0_startofpacket -> rsp_xbar_mux_001:sink64_startofpacket
	wire  [102:0] rsp_xbar_demux_064_src0_data;                                                                     // rsp_xbar_demux_064:src0_data -> rsp_xbar_mux_001:sink64_data
	wire   [98:0] rsp_xbar_demux_064_src0_channel;                                                                  // rsp_xbar_demux_064:src0_channel -> rsp_xbar_mux_001:sink64_channel
	wire          rsp_xbar_demux_064_src0_ready;                                                                    // rsp_xbar_mux_001:sink64_ready -> rsp_xbar_demux_064:src0_ready
	wire          rsp_xbar_demux_065_src0_endofpacket;                                                              // rsp_xbar_demux_065:src0_endofpacket -> rsp_xbar_mux_001:sink65_endofpacket
	wire          rsp_xbar_demux_065_src0_valid;                                                                    // rsp_xbar_demux_065:src0_valid -> rsp_xbar_mux_001:sink65_valid
	wire          rsp_xbar_demux_065_src0_startofpacket;                                                            // rsp_xbar_demux_065:src0_startofpacket -> rsp_xbar_mux_001:sink65_startofpacket
	wire  [102:0] rsp_xbar_demux_065_src0_data;                                                                     // rsp_xbar_demux_065:src0_data -> rsp_xbar_mux_001:sink65_data
	wire   [98:0] rsp_xbar_demux_065_src0_channel;                                                                  // rsp_xbar_demux_065:src0_channel -> rsp_xbar_mux_001:sink65_channel
	wire          rsp_xbar_demux_065_src0_ready;                                                                    // rsp_xbar_mux_001:sink65_ready -> rsp_xbar_demux_065:src0_ready
	wire          rsp_xbar_demux_066_src0_endofpacket;                                                              // rsp_xbar_demux_066:src0_endofpacket -> rsp_xbar_mux_001:sink66_endofpacket
	wire          rsp_xbar_demux_066_src0_valid;                                                                    // rsp_xbar_demux_066:src0_valid -> rsp_xbar_mux_001:sink66_valid
	wire          rsp_xbar_demux_066_src0_startofpacket;                                                            // rsp_xbar_demux_066:src0_startofpacket -> rsp_xbar_mux_001:sink66_startofpacket
	wire  [102:0] rsp_xbar_demux_066_src0_data;                                                                     // rsp_xbar_demux_066:src0_data -> rsp_xbar_mux_001:sink66_data
	wire   [98:0] rsp_xbar_demux_066_src0_channel;                                                                  // rsp_xbar_demux_066:src0_channel -> rsp_xbar_mux_001:sink66_channel
	wire          rsp_xbar_demux_066_src0_ready;                                                                    // rsp_xbar_mux_001:sink66_ready -> rsp_xbar_demux_066:src0_ready
	wire          rsp_xbar_demux_067_src0_endofpacket;                                                              // rsp_xbar_demux_067:src0_endofpacket -> rsp_xbar_mux_001:sink67_endofpacket
	wire          rsp_xbar_demux_067_src0_valid;                                                                    // rsp_xbar_demux_067:src0_valid -> rsp_xbar_mux_001:sink67_valid
	wire          rsp_xbar_demux_067_src0_startofpacket;                                                            // rsp_xbar_demux_067:src0_startofpacket -> rsp_xbar_mux_001:sink67_startofpacket
	wire  [102:0] rsp_xbar_demux_067_src0_data;                                                                     // rsp_xbar_demux_067:src0_data -> rsp_xbar_mux_001:sink67_data
	wire   [98:0] rsp_xbar_demux_067_src0_channel;                                                                  // rsp_xbar_demux_067:src0_channel -> rsp_xbar_mux_001:sink67_channel
	wire          rsp_xbar_demux_067_src0_ready;                                                                    // rsp_xbar_mux_001:sink67_ready -> rsp_xbar_demux_067:src0_ready
	wire          rsp_xbar_demux_068_src0_endofpacket;                                                              // rsp_xbar_demux_068:src0_endofpacket -> rsp_xbar_mux_001:sink68_endofpacket
	wire          rsp_xbar_demux_068_src0_valid;                                                                    // rsp_xbar_demux_068:src0_valid -> rsp_xbar_mux_001:sink68_valid
	wire          rsp_xbar_demux_068_src0_startofpacket;                                                            // rsp_xbar_demux_068:src0_startofpacket -> rsp_xbar_mux_001:sink68_startofpacket
	wire  [102:0] rsp_xbar_demux_068_src0_data;                                                                     // rsp_xbar_demux_068:src0_data -> rsp_xbar_mux_001:sink68_data
	wire   [98:0] rsp_xbar_demux_068_src0_channel;                                                                  // rsp_xbar_demux_068:src0_channel -> rsp_xbar_mux_001:sink68_channel
	wire          rsp_xbar_demux_068_src0_ready;                                                                    // rsp_xbar_mux_001:sink68_ready -> rsp_xbar_demux_068:src0_ready
	wire          rsp_xbar_demux_069_src0_endofpacket;                                                              // rsp_xbar_demux_069:src0_endofpacket -> rsp_xbar_mux_001:sink69_endofpacket
	wire          rsp_xbar_demux_069_src0_valid;                                                                    // rsp_xbar_demux_069:src0_valid -> rsp_xbar_mux_001:sink69_valid
	wire          rsp_xbar_demux_069_src0_startofpacket;                                                            // rsp_xbar_demux_069:src0_startofpacket -> rsp_xbar_mux_001:sink69_startofpacket
	wire  [102:0] rsp_xbar_demux_069_src0_data;                                                                     // rsp_xbar_demux_069:src0_data -> rsp_xbar_mux_001:sink69_data
	wire   [98:0] rsp_xbar_demux_069_src0_channel;                                                                  // rsp_xbar_demux_069:src0_channel -> rsp_xbar_mux_001:sink69_channel
	wire          rsp_xbar_demux_069_src0_ready;                                                                    // rsp_xbar_mux_001:sink69_ready -> rsp_xbar_demux_069:src0_ready
	wire          rsp_xbar_demux_070_src0_endofpacket;                                                              // rsp_xbar_demux_070:src0_endofpacket -> rsp_xbar_mux_001:sink70_endofpacket
	wire          rsp_xbar_demux_070_src0_valid;                                                                    // rsp_xbar_demux_070:src0_valid -> rsp_xbar_mux_001:sink70_valid
	wire          rsp_xbar_demux_070_src0_startofpacket;                                                            // rsp_xbar_demux_070:src0_startofpacket -> rsp_xbar_mux_001:sink70_startofpacket
	wire  [102:0] rsp_xbar_demux_070_src0_data;                                                                     // rsp_xbar_demux_070:src0_data -> rsp_xbar_mux_001:sink70_data
	wire   [98:0] rsp_xbar_demux_070_src0_channel;                                                                  // rsp_xbar_demux_070:src0_channel -> rsp_xbar_mux_001:sink70_channel
	wire          rsp_xbar_demux_070_src0_ready;                                                                    // rsp_xbar_mux_001:sink70_ready -> rsp_xbar_demux_070:src0_ready
	wire          rsp_xbar_demux_071_src0_endofpacket;                                                              // rsp_xbar_demux_071:src0_endofpacket -> rsp_xbar_mux_001:sink71_endofpacket
	wire          rsp_xbar_demux_071_src0_valid;                                                                    // rsp_xbar_demux_071:src0_valid -> rsp_xbar_mux_001:sink71_valid
	wire          rsp_xbar_demux_071_src0_startofpacket;                                                            // rsp_xbar_demux_071:src0_startofpacket -> rsp_xbar_mux_001:sink71_startofpacket
	wire  [102:0] rsp_xbar_demux_071_src0_data;                                                                     // rsp_xbar_demux_071:src0_data -> rsp_xbar_mux_001:sink71_data
	wire   [98:0] rsp_xbar_demux_071_src0_channel;                                                                  // rsp_xbar_demux_071:src0_channel -> rsp_xbar_mux_001:sink71_channel
	wire          rsp_xbar_demux_071_src0_ready;                                                                    // rsp_xbar_mux_001:sink71_ready -> rsp_xbar_demux_071:src0_ready
	wire          rsp_xbar_demux_072_src0_endofpacket;                                                              // rsp_xbar_demux_072:src0_endofpacket -> rsp_xbar_mux_001:sink72_endofpacket
	wire          rsp_xbar_demux_072_src0_valid;                                                                    // rsp_xbar_demux_072:src0_valid -> rsp_xbar_mux_001:sink72_valid
	wire          rsp_xbar_demux_072_src0_startofpacket;                                                            // rsp_xbar_demux_072:src0_startofpacket -> rsp_xbar_mux_001:sink72_startofpacket
	wire  [102:0] rsp_xbar_demux_072_src0_data;                                                                     // rsp_xbar_demux_072:src0_data -> rsp_xbar_mux_001:sink72_data
	wire   [98:0] rsp_xbar_demux_072_src0_channel;                                                                  // rsp_xbar_demux_072:src0_channel -> rsp_xbar_mux_001:sink72_channel
	wire          rsp_xbar_demux_072_src0_ready;                                                                    // rsp_xbar_mux_001:sink72_ready -> rsp_xbar_demux_072:src0_ready
	wire          rsp_xbar_demux_073_src0_endofpacket;                                                              // rsp_xbar_demux_073:src0_endofpacket -> rsp_xbar_mux_001:sink73_endofpacket
	wire          rsp_xbar_demux_073_src0_valid;                                                                    // rsp_xbar_demux_073:src0_valid -> rsp_xbar_mux_001:sink73_valid
	wire          rsp_xbar_demux_073_src0_startofpacket;                                                            // rsp_xbar_demux_073:src0_startofpacket -> rsp_xbar_mux_001:sink73_startofpacket
	wire  [102:0] rsp_xbar_demux_073_src0_data;                                                                     // rsp_xbar_demux_073:src0_data -> rsp_xbar_mux_001:sink73_data
	wire   [98:0] rsp_xbar_demux_073_src0_channel;                                                                  // rsp_xbar_demux_073:src0_channel -> rsp_xbar_mux_001:sink73_channel
	wire          rsp_xbar_demux_073_src0_ready;                                                                    // rsp_xbar_mux_001:sink73_ready -> rsp_xbar_demux_073:src0_ready
	wire          rsp_xbar_demux_074_src0_endofpacket;                                                              // rsp_xbar_demux_074:src0_endofpacket -> rsp_xbar_mux_001:sink74_endofpacket
	wire          rsp_xbar_demux_074_src0_valid;                                                                    // rsp_xbar_demux_074:src0_valid -> rsp_xbar_mux_001:sink74_valid
	wire          rsp_xbar_demux_074_src0_startofpacket;                                                            // rsp_xbar_demux_074:src0_startofpacket -> rsp_xbar_mux_001:sink74_startofpacket
	wire  [102:0] rsp_xbar_demux_074_src0_data;                                                                     // rsp_xbar_demux_074:src0_data -> rsp_xbar_mux_001:sink74_data
	wire   [98:0] rsp_xbar_demux_074_src0_channel;                                                                  // rsp_xbar_demux_074:src0_channel -> rsp_xbar_mux_001:sink74_channel
	wire          rsp_xbar_demux_074_src0_ready;                                                                    // rsp_xbar_mux_001:sink74_ready -> rsp_xbar_demux_074:src0_ready
	wire          rsp_xbar_demux_075_src0_endofpacket;                                                              // rsp_xbar_demux_075:src0_endofpacket -> rsp_xbar_mux_001:sink75_endofpacket
	wire          rsp_xbar_demux_075_src0_valid;                                                                    // rsp_xbar_demux_075:src0_valid -> rsp_xbar_mux_001:sink75_valid
	wire          rsp_xbar_demux_075_src0_startofpacket;                                                            // rsp_xbar_demux_075:src0_startofpacket -> rsp_xbar_mux_001:sink75_startofpacket
	wire  [102:0] rsp_xbar_demux_075_src0_data;                                                                     // rsp_xbar_demux_075:src0_data -> rsp_xbar_mux_001:sink75_data
	wire   [98:0] rsp_xbar_demux_075_src0_channel;                                                                  // rsp_xbar_demux_075:src0_channel -> rsp_xbar_mux_001:sink75_channel
	wire          rsp_xbar_demux_075_src0_ready;                                                                    // rsp_xbar_mux_001:sink75_ready -> rsp_xbar_demux_075:src0_ready
	wire          rsp_xbar_demux_076_src0_endofpacket;                                                              // rsp_xbar_demux_076:src0_endofpacket -> rsp_xbar_mux_001:sink76_endofpacket
	wire          rsp_xbar_demux_076_src0_valid;                                                                    // rsp_xbar_demux_076:src0_valid -> rsp_xbar_mux_001:sink76_valid
	wire          rsp_xbar_demux_076_src0_startofpacket;                                                            // rsp_xbar_demux_076:src0_startofpacket -> rsp_xbar_mux_001:sink76_startofpacket
	wire  [102:0] rsp_xbar_demux_076_src0_data;                                                                     // rsp_xbar_demux_076:src0_data -> rsp_xbar_mux_001:sink76_data
	wire   [98:0] rsp_xbar_demux_076_src0_channel;                                                                  // rsp_xbar_demux_076:src0_channel -> rsp_xbar_mux_001:sink76_channel
	wire          rsp_xbar_demux_076_src0_ready;                                                                    // rsp_xbar_mux_001:sink76_ready -> rsp_xbar_demux_076:src0_ready
	wire          rsp_xbar_demux_077_src0_endofpacket;                                                              // rsp_xbar_demux_077:src0_endofpacket -> rsp_xbar_mux_001:sink77_endofpacket
	wire          rsp_xbar_demux_077_src0_valid;                                                                    // rsp_xbar_demux_077:src0_valid -> rsp_xbar_mux_001:sink77_valid
	wire          rsp_xbar_demux_077_src0_startofpacket;                                                            // rsp_xbar_demux_077:src0_startofpacket -> rsp_xbar_mux_001:sink77_startofpacket
	wire  [102:0] rsp_xbar_demux_077_src0_data;                                                                     // rsp_xbar_demux_077:src0_data -> rsp_xbar_mux_001:sink77_data
	wire   [98:0] rsp_xbar_demux_077_src0_channel;                                                                  // rsp_xbar_demux_077:src0_channel -> rsp_xbar_mux_001:sink77_channel
	wire          rsp_xbar_demux_077_src0_ready;                                                                    // rsp_xbar_mux_001:sink77_ready -> rsp_xbar_demux_077:src0_ready
	wire          rsp_xbar_demux_078_src0_endofpacket;                                                              // rsp_xbar_demux_078:src0_endofpacket -> rsp_xbar_mux_001:sink78_endofpacket
	wire          rsp_xbar_demux_078_src0_valid;                                                                    // rsp_xbar_demux_078:src0_valid -> rsp_xbar_mux_001:sink78_valid
	wire          rsp_xbar_demux_078_src0_startofpacket;                                                            // rsp_xbar_demux_078:src0_startofpacket -> rsp_xbar_mux_001:sink78_startofpacket
	wire  [102:0] rsp_xbar_demux_078_src0_data;                                                                     // rsp_xbar_demux_078:src0_data -> rsp_xbar_mux_001:sink78_data
	wire   [98:0] rsp_xbar_demux_078_src0_channel;                                                                  // rsp_xbar_demux_078:src0_channel -> rsp_xbar_mux_001:sink78_channel
	wire          rsp_xbar_demux_078_src0_ready;                                                                    // rsp_xbar_mux_001:sink78_ready -> rsp_xbar_demux_078:src0_ready
	wire          rsp_xbar_demux_079_src0_endofpacket;                                                              // rsp_xbar_demux_079:src0_endofpacket -> rsp_xbar_mux_001:sink79_endofpacket
	wire          rsp_xbar_demux_079_src0_valid;                                                                    // rsp_xbar_demux_079:src0_valid -> rsp_xbar_mux_001:sink79_valid
	wire          rsp_xbar_demux_079_src0_startofpacket;                                                            // rsp_xbar_demux_079:src0_startofpacket -> rsp_xbar_mux_001:sink79_startofpacket
	wire  [102:0] rsp_xbar_demux_079_src0_data;                                                                     // rsp_xbar_demux_079:src0_data -> rsp_xbar_mux_001:sink79_data
	wire   [98:0] rsp_xbar_demux_079_src0_channel;                                                                  // rsp_xbar_demux_079:src0_channel -> rsp_xbar_mux_001:sink79_channel
	wire          rsp_xbar_demux_079_src0_ready;                                                                    // rsp_xbar_mux_001:sink79_ready -> rsp_xbar_demux_079:src0_ready
	wire          rsp_xbar_demux_080_src0_endofpacket;                                                              // rsp_xbar_demux_080:src0_endofpacket -> rsp_xbar_mux_001:sink80_endofpacket
	wire          rsp_xbar_demux_080_src0_valid;                                                                    // rsp_xbar_demux_080:src0_valid -> rsp_xbar_mux_001:sink80_valid
	wire          rsp_xbar_demux_080_src0_startofpacket;                                                            // rsp_xbar_demux_080:src0_startofpacket -> rsp_xbar_mux_001:sink80_startofpacket
	wire  [102:0] rsp_xbar_demux_080_src0_data;                                                                     // rsp_xbar_demux_080:src0_data -> rsp_xbar_mux_001:sink80_data
	wire   [98:0] rsp_xbar_demux_080_src0_channel;                                                                  // rsp_xbar_demux_080:src0_channel -> rsp_xbar_mux_001:sink80_channel
	wire          rsp_xbar_demux_080_src0_ready;                                                                    // rsp_xbar_mux_001:sink80_ready -> rsp_xbar_demux_080:src0_ready
	wire          rsp_xbar_demux_081_src0_endofpacket;                                                              // rsp_xbar_demux_081:src0_endofpacket -> rsp_xbar_mux_001:sink81_endofpacket
	wire          rsp_xbar_demux_081_src0_valid;                                                                    // rsp_xbar_demux_081:src0_valid -> rsp_xbar_mux_001:sink81_valid
	wire          rsp_xbar_demux_081_src0_startofpacket;                                                            // rsp_xbar_demux_081:src0_startofpacket -> rsp_xbar_mux_001:sink81_startofpacket
	wire  [102:0] rsp_xbar_demux_081_src0_data;                                                                     // rsp_xbar_demux_081:src0_data -> rsp_xbar_mux_001:sink81_data
	wire   [98:0] rsp_xbar_demux_081_src0_channel;                                                                  // rsp_xbar_demux_081:src0_channel -> rsp_xbar_mux_001:sink81_channel
	wire          rsp_xbar_demux_081_src0_ready;                                                                    // rsp_xbar_mux_001:sink81_ready -> rsp_xbar_demux_081:src0_ready
	wire          rsp_xbar_demux_082_src0_endofpacket;                                                              // rsp_xbar_demux_082:src0_endofpacket -> rsp_xbar_mux_001:sink82_endofpacket
	wire          rsp_xbar_demux_082_src0_valid;                                                                    // rsp_xbar_demux_082:src0_valid -> rsp_xbar_mux_001:sink82_valid
	wire          rsp_xbar_demux_082_src0_startofpacket;                                                            // rsp_xbar_demux_082:src0_startofpacket -> rsp_xbar_mux_001:sink82_startofpacket
	wire  [102:0] rsp_xbar_demux_082_src0_data;                                                                     // rsp_xbar_demux_082:src0_data -> rsp_xbar_mux_001:sink82_data
	wire   [98:0] rsp_xbar_demux_082_src0_channel;                                                                  // rsp_xbar_demux_082:src0_channel -> rsp_xbar_mux_001:sink82_channel
	wire          rsp_xbar_demux_082_src0_ready;                                                                    // rsp_xbar_mux_001:sink82_ready -> rsp_xbar_demux_082:src0_ready
	wire          rsp_xbar_demux_083_src0_endofpacket;                                                              // rsp_xbar_demux_083:src0_endofpacket -> rsp_xbar_mux_001:sink83_endofpacket
	wire          rsp_xbar_demux_083_src0_valid;                                                                    // rsp_xbar_demux_083:src0_valid -> rsp_xbar_mux_001:sink83_valid
	wire          rsp_xbar_demux_083_src0_startofpacket;                                                            // rsp_xbar_demux_083:src0_startofpacket -> rsp_xbar_mux_001:sink83_startofpacket
	wire  [102:0] rsp_xbar_demux_083_src0_data;                                                                     // rsp_xbar_demux_083:src0_data -> rsp_xbar_mux_001:sink83_data
	wire   [98:0] rsp_xbar_demux_083_src0_channel;                                                                  // rsp_xbar_demux_083:src0_channel -> rsp_xbar_mux_001:sink83_channel
	wire          rsp_xbar_demux_083_src0_ready;                                                                    // rsp_xbar_mux_001:sink83_ready -> rsp_xbar_demux_083:src0_ready
	wire          rsp_xbar_demux_084_src0_endofpacket;                                                              // rsp_xbar_demux_084:src0_endofpacket -> rsp_xbar_mux_001:sink84_endofpacket
	wire          rsp_xbar_demux_084_src0_valid;                                                                    // rsp_xbar_demux_084:src0_valid -> rsp_xbar_mux_001:sink84_valid
	wire          rsp_xbar_demux_084_src0_startofpacket;                                                            // rsp_xbar_demux_084:src0_startofpacket -> rsp_xbar_mux_001:sink84_startofpacket
	wire  [102:0] rsp_xbar_demux_084_src0_data;                                                                     // rsp_xbar_demux_084:src0_data -> rsp_xbar_mux_001:sink84_data
	wire   [98:0] rsp_xbar_demux_084_src0_channel;                                                                  // rsp_xbar_demux_084:src0_channel -> rsp_xbar_mux_001:sink84_channel
	wire          rsp_xbar_demux_084_src0_ready;                                                                    // rsp_xbar_mux_001:sink84_ready -> rsp_xbar_demux_084:src0_ready
	wire          rsp_xbar_demux_085_src0_endofpacket;                                                              // rsp_xbar_demux_085:src0_endofpacket -> rsp_xbar_mux_001:sink85_endofpacket
	wire          rsp_xbar_demux_085_src0_valid;                                                                    // rsp_xbar_demux_085:src0_valid -> rsp_xbar_mux_001:sink85_valid
	wire          rsp_xbar_demux_085_src0_startofpacket;                                                            // rsp_xbar_demux_085:src0_startofpacket -> rsp_xbar_mux_001:sink85_startofpacket
	wire  [102:0] rsp_xbar_demux_085_src0_data;                                                                     // rsp_xbar_demux_085:src0_data -> rsp_xbar_mux_001:sink85_data
	wire   [98:0] rsp_xbar_demux_085_src0_channel;                                                                  // rsp_xbar_demux_085:src0_channel -> rsp_xbar_mux_001:sink85_channel
	wire          rsp_xbar_demux_085_src0_ready;                                                                    // rsp_xbar_mux_001:sink85_ready -> rsp_xbar_demux_085:src0_ready
	wire          rsp_xbar_demux_086_src0_endofpacket;                                                              // rsp_xbar_demux_086:src0_endofpacket -> rsp_xbar_mux_001:sink86_endofpacket
	wire          rsp_xbar_demux_086_src0_valid;                                                                    // rsp_xbar_demux_086:src0_valid -> rsp_xbar_mux_001:sink86_valid
	wire          rsp_xbar_demux_086_src0_startofpacket;                                                            // rsp_xbar_demux_086:src0_startofpacket -> rsp_xbar_mux_001:sink86_startofpacket
	wire  [102:0] rsp_xbar_demux_086_src0_data;                                                                     // rsp_xbar_demux_086:src0_data -> rsp_xbar_mux_001:sink86_data
	wire   [98:0] rsp_xbar_demux_086_src0_channel;                                                                  // rsp_xbar_demux_086:src0_channel -> rsp_xbar_mux_001:sink86_channel
	wire          rsp_xbar_demux_086_src0_ready;                                                                    // rsp_xbar_mux_001:sink86_ready -> rsp_xbar_demux_086:src0_ready
	wire          rsp_xbar_demux_087_src0_endofpacket;                                                              // rsp_xbar_demux_087:src0_endofpacket -> rsp_xbar_mux_001:sink87_endofpacket
	wire          rsp_xbar_demux_087_src0_valid;                                                                    // rsp_xbar_demux_087:src0_valid -> rsp_xbar_mux_001:sink87_valid
	wire          rsp_xbar_demux_087_src0_startofpacket;                                                            // rsp_xbar_demux_087:src0_startofpacket -> rsp_xbar_mux_001:sink87_startofpacket
	wire  [102:0] rsp_xbar_demux_087_src0_data;                                                                     // rsp_xbar_demux_087:src0_data -> rsp_xbar_mux_001:sink87_data
	wire   [98:0] rsp_xbar_demux_087_src0_channel;                                                                  // rsp_xbar_demux_087:src0_channel -> rsp_xbar_mux_001:sink87_channel
	wire          rsp_xbar_demux_087_src0_ready;                                                                    // rsp_xbar_mux_001:sink87_ready -> rsp_xbar_demux_087:src0_ready
	wire          rsp_xbar_demux_088_src0_endofpacket;                                                              // rsp_xbar_demux_088:src0_endofpacket -> rsp_xbar_mux_001:sink88_endofpacket
	wire          rsp_xbar_demux_088_src0_valid;                                                                    // rsp_xbar_demux_088:src0_valid -> rsp_xbar_mux_001:sink88_valid
	wire          rsp_xbar_demux_088_src0_startofpacket;                                                            // rsp_xbar_demux_088:src0_startofpacket -> rsp_xbar_mux_001:sink88_startofpacket
	wire  [102:0] rsp_xbar_demux_088_src0_data;                                                                     // rsp_xbar_demux_088:src0_data -> rsp_xbar_mux_001:sink88_data
	wire   [98:0] rsp_xbar_demux_088_src0_channel;                                                                  // rsp_xbar_demux_088:src0_channel -> rsp_xbar_mux_001:sink88_channel
	wire          rsp_xbar_demux_088_src0_ready;                                                                    // rsp_xbar_mux_001:sink88_ready -> rsp_xbar_demux_088:src0_ready
	wire          rsp_xbar_demux_089_src0_endofpacket;                                                              // rsp_xbar_demux_089:src0_endofpacket -> rsp_xbar_mux_001:sink89_endofpacket
	wire          rsp_xbar_demux_089_src0_valid;                                                                    // rsp_xbar_demux_089:src0_valid -> rsp_xbar_mux_001:sink89_valid
	wire          rsp_xbar_demux_089_src0_startofpacket;                                                            // rsp_xbar_demux_089:src0_startofpacket -> rsp_xbar_mux_001:sink89_startofpacket
	wire  [102:0] rsp_xbar_demux_089_src0_data;                                                                     // rsp_xbar_demux_089:src0_data -> rsp_xbar_mux_001:sink89_data
	wire   [98:0] rsp_xbar_demux_089_src0_channel;                                                                  // rsp_xbar_demux_089:src0_channel -> rsp_xbar_mux_001:sink89_channel
	wire          rsp_xbar_demux_089_src0_ready;                                                                    // rsp_xbar_mux_001:sink89_ready -> rsp_xbar_demux_089:src0_ready
	wire          rsp_xbar_demux_090_src0_endofpacket;                                                              // rsp_xbar_demux_090:src0_endofpacket -> rsp_xbar_mux_001:sink90_endofpacket
	wire          rsp_xbar_demux_090_src0_valid;                                                                    // rsp_xbar_demux_090:src0_valid -> rsp_xbar_mux_001:sink90_valid
	wire          rsp_xbar_demux_090_src0_startofpacket;                                                            // rsp_xbar_demux_090:src0_startofpacket -> rsp_xbar_mux_001:sink90_startofpacket
	wire  [102:0] rsp_xbar_demux_090_src0_data;                                                                     // rsp_xbar_demux_090:src0_data -> rsp_xbar_mux_001:sink90_data
	wire   [98:0] rsp_xbar_demux_090_src0_channel;                                                                  // rsp_xbar_demux_090:src0_channel -> rsp_xbar_mux_001:sink90_channel
	wire          rsp_xbar_demux_090_src0_ready;                                                                    // rsp_xbar_mux_001:sink90_ready -> rsp_xbar_demux_090:src0_ready
	wire          rsp_xbar_demux_091_src0_endofpacket;                                                              // rsp_xbar_demux_091:src0_endofpacket -> rsp_xbar_mux_001:sink91_endofpacket
	wire          rsp_xbar_demux_091_src0_valid;                                                                    // rsp_xbar_demux_091:src0_valid -> rsp_xbar_mux_001:sink91_valid
	wire          rsp_xbar_demux_091_src0_startofpacket;                                                            // rsp_xbar_demux_091:src0_startofpacket -> rsp_xbar_mux_001:sink91_startofpacket
	wire  [102:0] rsp_xbar_demux_091_src0_data;                                                                     // rsp_xbar_demux_091:src0_data -> rsp_xbar_mux_001:sink91_data
	wire   [98:0] rsp_xbar_demux_091_src0_channel;                                                                  // rsp_xbar_demux_091:src0_channel -> rsp_xbar_mux_001:sink91_channel
	wire          rsp_xbar_demux_091_src0_ready;                                                                    // rsp_xbar_mux_001:sink91_ready -> rsp_xbar_demux_091:src0_ready
	wire          rsp_xbar_demux_092_src0_endofpacket;                                                              // rsp_xbar_demux_092:src0_endofpacket -> rsp_xbar_mux_001:sink92_endofpacket
	wire          rsp_xbar_demux_092_src0_valid;                                                                    // rsp_xbar_demux_092:src0_valid -> rsp_xbar_mux_001:sink92_valid
	wire          rsp_xbar_demux_092_src0_startofpacket;                                                            // rsp_xbar_demux_092:src0_startofpacket -> rsp_xbar_mux_001:sink92_startofpacket
	wire  [102:0] rsp_xbar_demux_092_src0_data;                                                                     // rsp_xbar_demux_092:src0_data -> rsp_xbar_mux_001:sink92_data
	wire   [98:0] rsp_xbar_demux_092_src0_channel;                                                                  // rsp_xbar_demux_092:src0_channel -> rsp_xbar_mux_001:sink92_channel
	wire          rsp_xbar_demux_092_src0_ready;                                                                    // rsp_xbar_mux_001:sink92_ready -> rsp_xbar_demux_092:src0_ready
	wire          rsp_xbar_demux_093_src0_endofpacket;                                                              // rsp_xbar_demux_093:src0_endofpacket -> rsp_xbar_mux_001:sink93_endofpacket
	wire          rsp_xbar_demux_093_src0_valid;                                                                    // rsp_xbar_demux_093:src0_valid -> rsp_xbar_mux_001:sink93_valid
	wire          rsp_xbar_demux_093_src0_startofpacket;                                                            // rsp_xbar_demux_093:src0_startofpacket -> rsp_xbar_mux_001:sink93_startofpacket
	wire  [102:0] rsp_xbar_demux_093_src0_data;                                                                     // rsp_xbar_demux_093:src0_data -> rsp_xbar_mux_001:sink93_data
	wire   [98:0] rsp_xbar_demux_093_src0_channel;                                                                  // rsp_xbar_demux_093:src0_channel -> rsp_xbar_mux_001:sink93_channel
	wire          rsp_xbar_demux_093_src0_ready;                                                                    // rsp_xbar_mux_001:sink93_ready -> rsp_xbar_demux_093:src0_ready
	wire          rsp_xbar_demux_094_src0_endofpacket;                                                              // rsp_xbar_demux_094:src0_endofpacket -> rsp_xbar_mux_001:sink94_endofpacket
	wire          rsp_xbar_demux_094_src0_valid;                                                                    // rsp_xbar_demux_094:src0_valid -> rsp_xbar_mux_001:sink94_valid
	wire          rsp_xbar_demux_094_src0_startofpacket;                                                            // rsp_xbar_demux_094:src0_startofpacket -> rsp_xbar_mux_001:sink94_startofpacket
	wire  [102:0] rsp_xbar_demux_094_src0_data;                                                                     // rsp_xbar_demux_094:src0_data -> rsp_xbar_mux_001:sink94_data
	wire   [98:0] rsp_xbar_demux_094_src0_channel;                                                                  // rsp_xbar_demux_094:src0_channel -> rsp_xbar_mux_001:sink94_channel
	wire          rsp_xbar_demux_094_src0_ready;                                                                    // rsp_xbar_mux_001:sink94_ready -> rsp_xbar_demux_094:src0_ready
	wire          rsp_xbar_demux_095_src0_endofpacket;                                                              // rsp_xbar_demux_095:src0_endofpacket -> rsp_xbar_mux_001:sink95_endofpacket
	wire          rsp_xbar_demux_095_src0_valid;                                                                    // rsp_xbar_demux_095:src0_valid -> rsp_xbar_mux_001:sink95_valid
	wire          rsp_xbar_demux_095_src0_startofpacket;                                                            // rsp_xbar_demux_095:src0_startofpacket -> rsp_xbar_mux_001:sink95_startofpacket
	wire  [102:0] rsp_xbar_demux_095_src0_data;                                                                     // rsp_xbar_demux_095:src0_data -> rsp_xbar_mux_001:sink95_data
	wire   [98:0] rsp_xbar_demux_095_src0_channel;                                                                  // rsp_xbar_demux_095:src0_channel -> rsp_xbar_mux_001:sink95_channel
	wire          rsp_xbar_demux_095_src0_ready;                                                                    // rsp_xbar_mux_001:sink95_ready -> rsp_xbar_demux_095:src0_ready
	wire          rsp_xbar_demux_096_src0_endofpacket;                                                              // rsp_xbar_demux_096:src0_endofpacket -> rsp_xbar_mux_001:sink96_endofpacket
	wire          rsp_xbar_demux_096_src0_valid;                                                                    // rsp_xbar_demux_096:src0_valid -> rsp_xbar_mux_001:sink96_valid
	wire          rsp_xbar_demux_096_src0_startofpacket;                                                            // rsp_xbar_demux_096:src0_startofpacket -> rsp_xbar_mux_001:sink96_startofpacket
	wire  [102:0] rsp_xbar_demux_096_src0_data;                                                                     // rsp_xbar_demux_096:src0_data -> rsp_xbar_mux_001:sink96_data
	wire   [98:0] rsp_xbar_demux_096_src0_channel;                                                                  // rsp_xbar_demux_096:src0_channel -> rsp_xbar_mux_001:sink96_channel
	wire          rsp_xbar_demux_096_src0_ready;                                                                    // rsp_xbar_mux_001:sink96_ready -> rsp_xbar_demux_096:src0_ready
	wire          rsp_xbar_demux_097_src0_endofpacket;                                                              // rsp_xbar_demux_097:src0_endofpacket -> rsp_xbar_mux_001:sink97_endofpacket
	wire          rsp_xbar_demux_097_src0_valid;                                                                    // rsp_xbar_demux_097:src0_valid -> rsp_xbar_mux_001:sink97_valid
	wire          rsp_xbar_demux_097_src0_startofpacket;                                                            // rsp_xbar_demux_097:src0_startofpacket -> rsp_xbar_mux_001:sink97_startofpacket
	wire  [102:0] rsp_xbar_demux_097_src0_data;                                                                     // rsp_xbar_demux_097:src0_data -> rsp_xbar_mux_001:sink97_data
	wire   [98:0] rsp_xbar_demux_097_src0_channel;                                                                  // rsp_xbar_demux_097:src0_channel -> rsp_xbar_mux_001:sink97_channel
	wire          rsp_xbar_demux_097_src0_ready;                                                                    // rsp_xbar_mux_001:sink97_ready -> rsp_xbar_demux_097:src0_ready
	wire          rsp_xbar_demux_098_src0_endofpacket;                                                              // rsp_xbar_demux_098:src0_endofpacket -> rsp_xbar_mux_001:sink98_endofpacket
	wire          rsp_xbar_demux_098_src0_valid;                                                                    // rsp_xbar_demux_098:src0_valid -> rsp_xbar_mux_001:sink98_valid
	wire          rsp_xbar_demux_098_src0_startofpacket;                                                            // rsp_xbar_demux_098:src0_startofpacket -> rsp_xbar_mux_001:sink98_startofpacket
	wire  [102:0] rsp_xbar_demux_098_src0_data;                                                                     // rsp_xbar_demux_098:src0_data -> rsp_xbar_mux_001:sink98_data
	wire   [98:0] rsp_xbar_demux_098_src0_channel;                                                                  // rsp_xbar_demux_098:src0_channel -> rsp_xbar_mux_001:sink98_channel
	wire          rsp_xbar_demux_098_src0_ready;                                                                    // rsp_xbar_mux_001:sink98_ready -> rsp_xbar_demux_098:src0_ready
	wire          addr_router_src_endofpacket;                                                                      // addr_router:src_endofpacket -> cmd_xbar_demux:sink_endofpacket
	wire          addr_router_src_valid;                                                                            // addr_router:src_valid -> cmd_xbar_demux:sink_valid
	wire          addr_router_src_startofpacket;                                                                    // addr_router:src_startofpacket -> cmd_xbar_demux:sink_startofpacket
	wire  [102:0] addr_router_src_data;                                                                             // addr_router:src_data -> cmd_xbar_demux:sink_data
	wire   [98:0] addr_router_src_channel;                                                                          // addr_router:src_channel -> cmd_xbar_demux:sink_channel
	wire          addr_router_src_ready;                                                                            // cmd_xbar_demux:sink_ready -> addr_router:src_ready
	wire          rsp_xbar_mux_src_endofpacket;                                                                     // rsp_xbar_mux:src_endofpacket -> NIOS_CPU_instruction_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          rsp_xbar_mux_src_valid;                                                                           // rsp_xbar_mux:src_valid -> NIOS_CPU_instruction_master_translator_avalon_universal_master_0_agent:rp_valid
	wire          rsp_xbar_mux_src_startofpacket;                                                                   // rsp_xbar_mux:src_startofpacket -> NIOS_CPU_instruction_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [102:0] rsp_xbar_mux_src_data;                                                                            // rsp_xbar_mux:src_data -> NIOS_CPU_instruction_master_translator_avalon_universal_master_0_agent:rp_data
	wire   [98:0] rsp_xbar_mux_src_channel;                                                                         // rsp_xbar_mux:src_channel -> NIOS_CPU_instruction_master_translator_avalon_universal_master_0_agent:rp_channel
	wire          rsp_xbar_mux_src_ready;                                                                           // NIOS_CPU_instruction_master_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_mux:src_ready
	wire          addr_router_001_src_endofpacket;                                                                  // addr_router_001:src_endofpacket -> cmd_xbar_demux_001:sink_endofpacket
	wire          addr_router_001_src_valid;                                                                        // addr_router_001:src_valid -> cmd_xbar_demux_001:sink_valid
	wire          addr_router_001_src_startofpacket;                                                                // addr_router_001:src_startofpacket -> cmd_xbar_demux_001:sink_startofpacket
	wire  [102:0] addr_router_001_src_data;                                                                         // addr_router_001:src_data -> cmd_xbar_demux_001:sink_data
	wire   [98:0] addr_router_001_src_channel;                                                                      // addr_router_001:src_channel -> cmd_xbar_demux_001:sink_channel
	wire          addr_router_001_src_ready;                                                                        // cmd_xbar_demux_001:sink_ready -> addr_router_001:src_ready
	wire          rsp_xbar_mux_001_src_endofpacket;                                                                 // rsp_xbar_mux_001:src_endofpacket -> NIOS_CPU_data_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          rsp_xbar_mux_001_src_valid;                                                                       // rsp_xbar_mux_001:src_valid -> NIOS_CPU_data_master_translator_avalon_universal_master_0_agent:rp_valid
	wire          rsp_xbar_mux_001_src_startofpacket;                                                               // rsp_xbar_mux_001:src_startofpacket -> NIOS_CPU_data_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [102:0] rsp_xbar_mux_001_src_data;                                                                        // rsp_xbar_mux_001:src_data -> NIOS_CPU_data_master_translator_avalon_universal_master_0_agent:rp_data
	wire   [98:0] rsp_xbar_mux_001_src_channel;                                                                     // rsp_xbar_mux_001:src_channel -> NIOS_CPU_data_master_translator_avalon_universal_master_0_agent:rp_channel
	wire          rsp_xbar_mux_001_src_ready;                                                                       // NIOS_CPU_data_master_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_mux_001:src_ready
	wire          cmd_xbar_mux_src_endofpacket;                                                                     // cmd_xbar_mux:src_endofpacket -> NIOS_CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_mux_src_valid;                                                                           // cmd_xbar_mux:src_valid -> NIOS_CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_mux_src_startofpacket;                                                                   // cmd_xbar_mux:src_startofpacket -> NIOS_CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] cmd_xbar_mux_src_data;                                                                            // cmd_xbar_mux:src_data -> NIOS_CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_data
	wire   [98:0] cmd_xbar_mux_src_channel;                                                                         // cmd_xbar_mux:src_channel -> NIOS_CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_mux_src_ready;                                                                           // NIOS_CPU_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux:src_ready
	wire          id_router_src_endofpacket;                                                                        // id_router:src_endofpacket -> rsp_xbar_demux:sink_endofpacket
	wire          id_router_src_valid;                                                                              // id_router:src_valid -> rsp_xbar_demux:sink_valid
	wire          id_router_src_startofpacket;                                                                      // id_router:src_startofpacket -> rsp_xbar_demux:sink_startofpacket
	wire  [102:0] id_router_src_data;                                                                               // id_router:src_data -> rsp_xbar_demux:sink_data
	wire   [98:0] id_router_src_channel;                                                                            // id_router:src_channel -> rsp_xbar_demux:sink_channel
	wire          id_router_src_ready;                                                                              // rsp_xbar_demux:sink_ready -> id_router:src_ready
	wire          cmd_xbar_mux_001_src_endofpacket;                                                                 // cmd_xbar_mux_001:src_endofpacket -> RAM_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_mux_001_src_valid;                                                                       // cmd_xbar_mux_001:src_valid -> RAM_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_mux_001_src_startofpacket;                                                               // cmd_xbar_mux_001:src_startofpacket -> RAM_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] cmd_xbar_mux_001_src_data;                                                                        // cmd_xbar_mux_001:src_data -> RAM_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [98:0] cmd_xbar_mux_001_src_channel;                                                                     // cmd_xbar_mux_001:src_channel -> RAM_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_mux_001_src_ready;                                                                       // RAM_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_001:src_ready
	wire          id_router_001_src_endofpacket;                                                                    // id_router_001:src_endofpacket -> rsp_xbar_demux_001:sink_endofpacket
	wire          id_router_001_src_valid;                                                                          // id_router_001:src_valid -> rsp_xbar_demux_001:sink_valid
	wire          id_router_001_src_startofpacket;                                                                  // id_router_001:src_startofpacket -> rsp_xbar_demux_001:sink_startofpacket
	wire  [102:0] id_router_001_src_data;                                                                           // id_router_001:src_data -> rsp_xbar_demux_001:sink_data
	wire   [98:0] id_router_001_src_channel;                                                                        // id_router_001:src_channel -> rsp_xbar_demux_001:sink_channel
	wire          id_router_001_src_ready;                                                                          // rsp_xbar_demux_001:sink_ready -> id_router_001:src_ready
	wire          cmd_xbar_mux_002_src_endofpacket;                                                                 // cmd_xbar_mux_002:src_endofpacket -> SSRAM_uas_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_mux_002_src_valid;                                                                       // cmd_xbar_mux_002:src_valid -> SSRAM_uas_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_mux_002_src_startofpacket;                                                               // cmd_xbar_mux_002:src_startofpacket -> SSRAM_uas_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] cmd_xbar_mux_002_src_data;                                                                        // cmd_xbar_mux_002:src_data -> SSRAM_uas_translator_avalon_universal_slave_0_agent:cp_data
	wire   [98:0] cmd_xbar_mux_002_src_channel;                                                                     // cmd_xbar_mux_002:src_channel -> SSRAM_uas_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_mux_002_src_ready;                                                                       // SSRAM_uas_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_002:src_ready
	wire          id_router_002_src_endofpacket;                                                                    // id_router_002:src_endofpacket -> rsp_xbar_demux_002:sink_endofpacket
	wire          id_router_002_src_valid;                                                                          // id_router_002:src_valid -> rsp_xbar_demux_002:sink_valid
	wire          id_router_002_src_startofpacket;                                                                  // id_router_002:src_startofpacket -> rsp_xbar_demux_002:sink_startofpacket
	wire  [102:0] id_router_002_src_data;                                                                           // id_router_002:src_data -> rsp_xbar_demux_002:sink_data
	wire   [98:0] id_router_002_src_channel;                                                                        // id_router_002:src_channel -> rsp_xbar_demux_002:sink_channel
	wire          id_router_002_src_ready;                                                                          // rsp_xbar_demux_002:sink_ready -> id_router_002:src_ready
	wire          cmd_xbar_demux_001_src3_ready;                                                                    // JTAG_UART_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src3_ready
	wire          id_router_003_src_endofpacket;                                                                    // id_router_003:src_endofpacket -> rsp_xbar_demux_003:sink_endofpacket
	wire          id_router_003_src_valid;                                                                          // id_router_003:src_valid -> rsp_xbar_demux_003:sink_valid
	wire          id_router_003_src_startofpacket;                                                                  // id_router_003:src_startofpacket -> rsp_xbar_demux_003:sink_startofpacket
	wire  [102:0] id_router_003_src_data;                                                                           // id_router_003:src_data -> rsp_xbar_demux_003:sink_data
	wire   [98:0] id_router_003_src_channel;                                                                        // id_router_003:src_channel -> rsp_xbar_demux_003:sink_channel
	wire          id_router_003_src_ready;                                                                          // rsp_xbar_demux_003:sink_ready -> id_router_003:src_ready
	wire          cmd_xbar_demux_001_src4_ready;                                                                    // LCD_control_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src4_ready
	wire          id_router_004_src_endofpacket;                                                                    // id_router_004:src_endofpacket -> rsp_xbar_demux_004:sink_endofpacket
	wire          id_router_004_src_valid;                                                                          // id_router_004:src_valid -> rsp_xbar_demux_004:sink_valid
	wire          id_router_004_src_startofpacket;                                                                  // id_router_004:src_startofpacket -> rsp_xbar_demux_004:sink_startofpacket
	wire  [102:0] id_router_004_src_data;                                                                           // id_router_004:src_data -> rsp_xbar_demux_004:sink_data
	wire   [98:0] id_router_004_src_channel;                                                                        // id_router_004:src_channel -> rsp_xbar_demux_004:sink_channel
	wire          id_router_004_src_ready;                                                                          // rsp_xbar_demux_004:sink_ready -> id_router_004:src_ready
	wire          cmd_xbar_demux_001_src5_ready;                                                                    // ADC_ON_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src5_ready
	wire          id_router_005_src_endofpacket;                                                                    // id_router_005:src_endofpacket -> rsp_xbar_demux_005:sink_endofpacket
	wire          id_router_005_src_valid;                                                                          // id_router_005:src_valid -> rsp_xbar_demux_005:sink_valid
	wire          id_router_005_src_startofpacket;                                                                  // id_router_005:src_startofpacket -> rsp_xbar_demux_005:sink_startofpacket
	wire  [102:0] id_router_005_src_data;                                                                           // id_router_005:src_data -> rsp_xbar_demux_005:sink_data
	wire   [98:0] id_router_005_src_channel;                                                                        // id_router_005:src_channel -> rsp_xbar_demux_005:sink_channel
	wire          id_router_005_src_ready;                                                                          // rsp_xbar_demux_005:sink_ready -> id_router_005:src_ready
	wire          cmd_xbar_demux_001_src6_ready;                                                                    // FIFO_ADC_DATA_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src6_ready
	wire          id_router_006_src_endofpacket;                                                                    // id_router_006:src_endofpacket -> rsp_xbar_demux_006:sink_endofpacket
	wire          id_router_006_src_valid;                                                                          // id_router_006:src_valid -> rsp_xbar_demux_006:sink_valid
	wire          id_router_006_src_startofpacket;                                                                  // id_router_006:src_startofpacket -> rsp_xbar_demux_006:sink_startofpacket
	wire  [102:0] id_router_006_src_data;                                                                           // id_router_006:src_data -> rsp_xbar_demux_006:sink_data
	wire   [98:0] id_router_006_src_channel;                                                                        // id_router_006:src_channel -> rsp_xbar_demux_006:sink_channel
	wire          id_router_006_src_ready;                                                                          // rsp_xbar_demux_006:sink_ready -> id_router_006:src_ready
	wire          cmd_xbar_demux_001_src7_ready;                                                                    // FIFO_ADC_DATA_VALID_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src7_ready
	wire          id_router_007_src_endofpacket;                                                                    // id_router_007:src_endofpacket -> rsp_xbar_demux_007:sink_endofpacket
	wire          id_router_007_src_valid;                                                                          // id_router_007:src_valid -> rsp_xbar_demux_007:sink_valid
	wire          id_router_007_src_startofpacket;                                                                  // id_router_007:src_startofpacket -> rsp_xbar_demux_007:sink_startofpacket
	wire  [102:0] id_router_007_src_data;                                                                           // id_router_007:src_data -> rsp_xbar_demux_007:sink_data
	wire   [98:0] id_router_007_src_channel;                                                                        // id_router_007:src_channel -> rsp_xbar_demux_007:sink_channel
	wire          id_router_007_src_ready;                                                                          // rsp_xbar_demux_007:sink_ready -> id_router_007:src_ready
	wire          cmd_xbar_demux_001_src8_ready;                                                                    // FIFO_RST_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src8_ready
	wire          id_router_008_src_endofpacket;                                                                    // id_router_008:src_endofpacket -> rsp_xbar_demux_008:sink_endofpacket
	wire          id_router_008_src_valid;                                                                          // id_router_008:src_valid -> rsp_xbar_demux_008:sink_valid
	wire          id_router_008_src_startofpacket;                                                                  // id_router_008:src_startofpacket -> rsp_xbar_demux_008:sink_startofpacket
	wire  [102:0] id_router_008_src_data;                                                                           // id_router_008:src_data -> rsp_xbar_demux_008:sink_data
	wire   [98:0] id_router_008_src_channel;                                                                        // id_router_008:src_channel -> rsp_xbar_demux_008:sink_channel
	wire          id_router_008_src_ready;                                                                          // rsp_xbar_demux_008:sink_ready -> id_router_008:src_ready
	wire          cmd_xbar_demux_001_src9_ready;                                                                    // SUBTRACTOR_ON_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src9_ready
	wire          id_router_009_src_endofpacket;                                                                    // id_router_009:src_endofpacket -> rsp_xbar_demux_009:sink_endofpacket
	wire          id_router_009_src_valid;                                                                          // id_router_009:src_valid -> rsp_xbar_demux_009:sink_valid
	wire          id_router_009_src_startofpacket;                                                                  // id_router_009:src_startofpacket -> rsp_xbar_demux_009:sink_startofpacket
	wire  [102:0] id_router_009_src_data;                                                                           // id_router_009:src_data -> rsp_xbar_demux_009:sink_data
	wire   [98:0] id_router_009_src_channel;                                                                        // id_router_009:src_channel -> rsp_xbar_demux_009:sink_channel
	wire          id_router_009_src_ready;                                                                          // rsp_xbar_demux_009:sink_ready -> id_router_009:src_ready
	wire          cmd_xbar_demux_001_src10_ready;                                                                   // CH0_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src10_ready
	wire          id_router_010_src_endofpacket;                                                                    // id_router_010:src_endofpacket -> rsp_xbar_demux_010:sink_endofpacket
	wire          id_router_010_src_valid;                                                                          // id_router_010:src_valid -> rsp_xbar_demux_010:sink_valid
	wire          id_router_010_src_startofpacket;                                                                  // id_router_010:src_startofpacket -> rsp_xbar_demux_010:sink_startofpacket
	wire  [102:0] id_router_010_src_data;                                                                           // id_router_010:src_data -> rsp_xbar_demux_010:sink_data
	wire   [98:0] id_router_010_src_channel;                                                                        // id_router_010:src_channel -> rsp_xbar_demux_010:sink_channel
	wire          id_router_010_src_ready;                                                                          // rsp_xbar_demux_010:sink_ready -> id_router_010:src_ready
	wire          cmd_xbar_demux_001_src11_ready;                                                                   // DETECTOR_ON_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src11_ready
	wire          id_router_011_src_endofpacket;                                                                    // id_router_011:src_endofpacket -> rsp_xbar_demux_011:sink_endofpacket
	wire          id_router_011_src_valid;                                                                          // id_router_011:src_valid -> rsp_xbar_demux_011:sink_valid
	wire          id_router_011_src_startofpacket;                                                                  // id_router_011:src_startofpacket -> rsp_xbar_demux_011:sink_startofpacket
	wire  [102:0] id_router_011_src_data;                                                                           // id_router_011:src_data -> rsp_xbar_demux_011:sink_data
	wire   [98:0] id_router_011_src_channel;                                                                        // id_router_011:src_channel -> rsp_xbar_demux_011:sink_channel
	wire          id_router_011_src_ready;                                                                          // rsp_xbar_demux_011:sink_ready -> id_router_011:src_ready
	wire          cmd_xbar_demux_001_src12_ready;                                                                   // MENU_DOWN_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src12_ready
	wire          id_router_012_src_endofpacket;                                                                    // id_router_012:src_endofpacket -> rsp_xbar_demux_012:sink_endofpacket
	wire          id_router_012_src_valid;                                                                          // id_router_012:src_valid -> rsp_xbar_demux_012:sink_valid
	wire          id_router_012_src_startofpacket;                                                                  // id_router_012:src_startofpacket -> rsp_xbar_demux_012:sink_startofpacket
	wire  [102:0] id_router_012_src_data;                                                                           // id_router_012:src_data -> rsp_xbar_demux_012:sink_data
	wire   [98:0] id_router_012_src_channel;                                                                        // id_router_012:src_channel -> rsp_xbar_demux_012:sink_channel
	wire          id_router_012_src_ready;                                                                          // rsp_xbar_demux_012:sink_ready -> id_router_012:src_ready
	wire          cmd_xbar_demux_001_src13_ready;                                                                   // MENU_UP_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src13_ready
	wire          id_router_013_src_endofpacket;                                                                    // id_router_013:src_endofpacket -> rsp_xbar_demux_013:sink_endofpacket
	wire          id_router_013_src_valid;                                                                          // id_router_013:src_valid -> rsp_xbar_demux_013:sink_valid
	wire          id_router_013_src_startofpacket;                                                                  // id_router_013:src_startofpacket -> rsp_xbar_demux_013:sink_startofpacket
	wire  [102:0] id_router_013_src_data;                                                                           // id_router_013:src_data -> rsp_xbar_demux_013:sink_data
	wire   [98:0] id_router_013_src_channel;                                                                        // id_router_013:src_channel -> rsp_xbar_demux_013:sink_channel
	wire          id_router_013_src_ready;                                                                          // rsp_xbar_demux_013:sink_ready -> id_router_013:src_ready
	wire          cmd_xbar_demux_001_src14_ready;                                                                   // MENU_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src14_ready
	wire          id_router_014_src_endofpacket;                                                                    // id_router_014:src_endofpacket -> rsp_xbar_demux_014:sink_endofpacket
	wire          id_router_014_src_valid;                                                                          // id_router_014:src_valid -> rsp_xbar_demux_014:sink_valid
	wire          id_router_014_src_startofpacket;                                                                  // id_router_014:src_startofpacket -> rsp_xbar_demux_014:sink_startofpacket
	wire  [102:0] id_router_014_src_data;                                                                           // id_router_014:src_data -> rsp_xbar_demux_014:sink_data
	wire   [98:0] id_router_014_src_channel;                                                                        // id_router_014:src_channel -> rsp_xbar_demux_014:sink_channel
	wire          id_router_014_src_ready;                                                                          // rsp_xbar_demux_014:sink_ready -> id_router_014:src_ready
	wire          cmd_xbar_demux_001_src15_ready;                                                                   // CH0_THRESH_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src15_ready
	wire          id_router_015_src_endofpacket;                                                                    // id_router_015:src_endofpacket -> rsp_xbar_demux_015:sink_endofpacket
	wire          id_router_015_src_valid;                                                                          // id_router_015:src_valid -> rsp_xbar_demux_015:sink_valid
	wire          id_router_015_src_startofpacket;                                                                  // id_router_015:src_startofpacket -> rsp_xbar_demux_015:sink_startofpacket
	wire  [102:0] id_router_015_src_data;                                                                           // id_router_015:src_data -> rsp_xbar_demux_015:sink_data
	wire   [98:0] id_router_015_src_channel;                                                                        // id_router_015:src_channel -> rsp_xbar_demux_015:sink_channel
	wire          id_router_015_src_ready;                                                                          // rsp_xbar_demux_015:sink_ready -> id_router_015:src_ready
	wire          cmd_xbar_demux_001_src16_ready;                                                                   // CH0_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src16_ready
	wire          id_router_016_src_endofpacket;                                                                    // id_router_016:src_endofpacket -> rsp_xbar_demux_016:sink_endofpacket
	wire          id_router_016_src_valid;                                                                          // id_router_016:src_valid -> rsp_xbar_demux_016:sink_valid
	wire          id_router_016_src_startofpacket;                                                                  // id_router_016:src_startofpacket -> rsp_xbar_demux_016:sink_startofpacket
	wire  [102:0] id_router_016_src_data;                                                                           // id_router_016:src_data -> rsp_xbar_demux_016:sink_data
	wire   [98:0] id_router_016_src_channel;                                                                        // id_router_016:src_channel -> rsp_xbar_demux_016:sink_channel
	wire          id_router_016_src_ready;                                                                          // rsp_xbar_demux_016:sink_ready -> id_router_016:src_ready
	wire          cmd_xbar_demux_001_src17_ready;                                                                   // CH0_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src17_ready
	wire          id_router_017_src_endofpacket;                                                                    // id_router_017:src_endofpacket -> rsp_xbar_demux_017:sink_endofpacket
	wire          id_router_017_src_valid;                                                                          // id_router_017:src_valid -> rsp_xbar_demux_017:sink_valid
	wire          id_router_017_src_startofpacket;                                                                  // id_router_017:src_startofpacket -> rsp_xbar_demux_017:sink_startofpacket
	wire  [102:0] id_router_017_src_data;                                                                           // id_router_017:src_data -> rsp_xbar_demux_017:sink_data
	wire   [98:0] id_router_017_src_channel;                                                                        // id_router_017:src_channel -> rsp_xbar_demux_017:sink_channel
	wire          id_router_017_src_ready;                                                                          // rsp_xbar_demux_017:sink_ready -> id_router_017:src_ready
	wire          cmd_xbar_demux_001_src18_ready;                                                                   // CH0_YN1_L_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src18_ready
	wire          id_router_018_src_endofpacket;                                                                    // id_router_018:src_endofpacket -> rsp_xbar_demux_018:sink_endofpacket
	wire          id_router_018_src_valid;                                                                          // id_router_018:src_valid -> rsp_xbar_demux_018:sink_valid
	wire          id_router_018_src_startofpacket;                                                                  // id_router_018:src_startofpacket -> rsp_xbar_demux_018:sink_startofpacket
	wire  [102:0] id_router_018_src_data;                                                                           // id_router_018:src_data -> rsp_xbar_demux_018:sink_data
	wire   [98:0] id_router_018_src_channel;                                                                        // id_router_018:src_channel -> rsp_xbar_demux_018:sink_channel
	wire          id_router_018_src_ready;                                                                          // rsp_xbar_demux_018:sink_ready -> id_router_018:src_ready
	wire          cmd_xbar_demux_001_src19_ready;                                                                   // CH0_YN1_ML_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src19_ready
	wire          id_router_019_src_endofpacket;                                                                    // id_router_019:src_endofpacket -> rsp_xbar_demux_019:sink_endofpacket
	wire          id_router_019_src_valid;                                                                          // id_router_019:src_valid -> rsp_xbar_demux_019:sink_valid
	wire          id_router_019_src_startofpacket;                                                                  // id_router_019:src_startofpacket -> rsp_xbar_demux_019:sink_startofpacket
	wire  [102:0] id_router_019_src_data;                                                                           // id_router_019:src_data -> rsp_xbar_demux_019:sink_data
	wire   [98:0] id_router_019_src_channel;                                                                        // id_router_019:src_channel -> rsp_xbar_demux_019:sink_channel
	wire          id_router_019_src_ready;                                                                          // rsp_xbar_demux_019:sink_ready -> id_router_019:src_ready
	wire          cmd_xbar_demux_001_src20_ready;                                                                   // CH0_YN1_MU_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src20_ready
	wire          id_router_020_src_endofpacket;                                                                    // id_router_020:src_endofpacket -> rsp_xbar_demux_020:sink_endofpacket
	wire          id_router_020_src_valid;                                                                          // id_router_020:src_valid -> rsp_xbar_demux_020:sink_valid
	wire          id_router_020_src_startofpacket;                                                                  // id_router_020:src_startofpacket -> rsp_xbar_demux_020:sink_startofpacket
	wire  [102:0] id_router_020_src_data;                                                                           // id_router_020:src_data -> rsp_xbar_demux_020:sink_data
	wire   [98:0] id_router_020_src_channel;                                                                        // id_router_020:src_channel -> rsp_xbar_demux_020:sink_channel
	wire          id_router_020_src_ready;                                                                          // rsp_xbar_demux_020:sink_ready -> id_router_020:src_ready
	wire          cmd_xbar_demux_001_src21_ready;                                                                   // CH0_YN1_U_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src21_ready
	wire          id_router_021_src_endofpacket;                                                                    // id_router_021:src_endofpacket -> rsp_xbar_demux_021:sink_endofpacket
	wire          id_router_021_src_valid;                                                                          // id_router_021:src_valid -> rsp_xbar_demux_021:sink_valid
	wire          id_router_021_src_startofpacket;                                                                  // id_router_021:src_startofpacket -> rsp_xbar_demux_021:sink_startofpacket
	wire  [102:0] id_router_021_src_data;                                                                           // id_router_021:src_data -> rsp_xbar_demux_021:sink_data
	wire   [98:0] id_router_021_src_channel;                                                                        // id_router_021:src_channel -> rsp_xbar_demux_021:sink_channel
	wire          id_router_021_src_ready;                                                                          // rsp_xbar_demux_021:sink_ready -> id_router_021:src_ready
	wire          cmd_xbar_demux_001_src22_ready;                                                                   // CH0_TIME_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src22_ready
	wire          id_router_022_src_endofpacket;                                                                    // id_router_022:src_endofpacket -> rsp_xbar_demux_022:sink_endofpacket
	wire          id_router_022_src_valid;                                                                          // id_router_022:src_valid -> rsp_xbar_demux_022:sink_valid
	wire          id_router_022_src_startofpacket;                                                                  // id_router_022:src_startofpacket -> rsp_xbar_demux_022:sink_startofpacket
	wire  [102:0] id_router_022_src_data;                                                                           // id_router_022:src_data -> rsp_xbar_demux_022:sink_data
	wire   [98:0] id_router_022_src_channel;                                                                        // id_router_022:src_channel -> rsp_xbar_demux_022:sink_channel
	wire          id_router_022_src_ready;                                                                          // rsp_xbar_demux_022:sink_ready -> id_router_022:src_ready
	wire          cmd_xbar_demux_001_src23_ready;                                                                   // CH0_YN2_MU_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src23_ready
	wire          id_router_023_src_endofpacket;                                                                    // id_router_023:src_endofpacket -> rsp_xbar_demux_023:sink_endofpacket
	wire          id_router_023_src_valid;                                                                          // id_router_023:src_valid -> rsp_xbar_demux_023:sink_valid
	wire          id_router_023_src_startofpacket;                                                                  // id_router_023:src_startofpacket -> rsp_xbar_demux_023:sink_startofpacket
	wire  [102:0] id_router_023_src_data;                                                                           // id_router_023:src_data -> rsp_xbar_demux_023:sink_data
	wire   [98:0] id_router_023_src_channel;                                                                        // id_router_023:src_channel -> rsp_xbar_demux_023:sink_channel
	wire          id_router_023_src_ready;                                                                          // rsp_xbar_demux_023:sink_ready -> id_router_023:src_ready
	wire          cmd_xbar_demux_001_src24_ready;                                                                   // CH0_YN2_ML_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src24_ready
	wire          id_router_024_src_endofpacket;                                                                    // id_router_024:src_endofpacket -> rsp_xbar_demux_024:sink_endofpacket
	wire          id_router_024_src_valid;                                                                          // id_router_024:src_valid -> rsp_xbar_demux_024:sink_valid
	wire          id_router_024_src_startofpacket;                                                                  // id_router_024:src_startofpacket -> rsp_xbar_demux_024:sink_startofpacket
	wire  [102:0] id_router_024_src_data;                                                                           // id_router_024:src_data -> rsp_xbar_demux_024:sink_data
	wire   [98:0] id_router_024_src_channel;                                                                        // id_router_024:src_channel -> rsp_xbar_demux_024:sink_channel
	wire          id_router_024_src_ready;                                                                          // rsp_xbar_demux_024:sink_ready -> id_router_024:src_ready
	wire          cmd_xbar_demux_001_src25_ready;                                                                   // CH0_YN2_U_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src25_ready
	wire          id_router_025_src_endofpacket;                                                                    // id_router_025:src_endofpacket -> rsp_xbar_demux_025:sink_endofpacket
	wire          id_router_025_src_valid;                                                                          // id_router_025:src_valid -> rsp_xbar_demux_025:sink_valid
	wire          id_router_025_src_startofpacket;                                                                  // id_router_025:src_startofpacket -> rsp_xbar_demux_025:sink_startofpacket
	wire  [102:0] id_router_025_src_data;                                                                           // id_router_025:src_data -> rsp_xbar_demux_025:sink_data
	wire   [98:0] id_router_025_src_channel;                                                                        // id_router_025:src_channel -> rsp_xbar_demux_025:sink_channel
	wire          id_router_025_src_ready;                                                                          // rsp_xbar_demux_025:sink_ready -> id_router_025:src_ready
	wire          cmd_xbar_demux_001_src26_ready;                                                                   // CH0_YN2_L_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src26_ready
	wire          id_router_026_src_endofpacket;                                                                    // id_router_026:src_endofpacket -> rsp_xbar_demux_026:sink_endofpacket
	wire          id_router_026_src_valid;                                                                          // id_router_026:src_valid -> rsp_xbar_demux_026:sink_valid
	wire          id_router_026_src_startofpacket;                                                                  // id_router_026:src_startofpacket -> rsp_xbar_demux_026:sink_startofpacket
	wire  [102:0] id_router_026_src_data;                                                                           // id_router_026:src_data -> rsp_xbar_demux_026:sink_data
	wire   [98:0] id_router_026_src_channel;                                                                        // id_router_026:src_channel -> rsp_xbar_demux_026:sink_channel
	wire          id_router_026_src_ready;                                                                          // rsp_xbar_demux_026:sink_ready -> id_router_026:src_ready
	wire          cmd_xbar_demux_001_src27_ready;                                                                   // CH0_YN3_L_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src27_ready
	wire          id_router_027_src_endofpacket;                                                                    // id_router_027:src_endofpacket -> rsp_xbar_demux_027:sink_endofpacket
	wire          id_router_027_src_valid;                                                                          // id_router_027:src_valid -> rsp_xbar_demux_027:sink_valid
	wire          id_router_027_src_startofpacket;                                                                  // id_router_027:src_startofpacket -> rsp_xbar_demux_027:sink_startofpacket
	wire  [102:0] id_router_027_src_data;                                                                           // id_router_027:src_data -> rsp_xbar_demux_027:sink_data
	wire   [98:0] id_router_027_src_channel;                                                                        // id_router_027:src_channel -> rsp_xbar_demux_027:sink_channel
	wire          id_router_027_src_ready;                                                                          // rsp_xbar_demux_027:sink_ready -> id_router_027:src_ready
	wire          cmd_xbar_demux_001_src28_ready;                                                                   // CH0_YN3_ML_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src28_ready
	wire          id_router_028_src_endofpacket;                                                                    // id_router_028:src_endofpacket -> rsp_xbar_demux_028:sink_endofpacket
	wire          id_router_028_src_valid;                                                                          // id_router_028:src_valid -> rsp_xbar_demux_028:sink_valid
	wire          id_router_028_src_startofpacket;                                                                  // id_router_028:src_startofpacket -> rsp_xbar_demux_028:sink_startofpacket
	wire  [102:0] id_router_028_src_data;                                                                           // id_router_028:src_data -> rsp_xbar_demux_028:sink_data
	wire   [98:0] id_router_028_src_channel;                                                                        // id_router_028:src_channel -> rsp_xbar_demux_028:sink_channel
	wire          id_router_028_src_ready;                                                                          // rsp_xbar_demux_028:sink_ready -> id_router_028:src_ready
	wire          cmd_xbar_demux_001_src29_ready;                                                                   // CH0_YN3_MU_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src29_ready
	wire          id_router_029_src_endofpacket;                                                                    // id_router_029:src_endofpacket -> rsp_xbar_demux_029:sink_endofpacket
	wire          id_router_029_src_valid;                                                                          // id_router_029:src_valid -> rsp_xbar_demux_029:sink_valid
	wire          id_router_029_src_startofpacket;                                                                  // id_router_029:src_startofpacket -> rsp_xbar_demux_029:sink_startofpacket
	wire  [102:0] id_router_029_src_data;                                                                           // id_router_029:src_data -> rsp_xbar_demux_029:sink_data
	wire   [98:0] id_router_029_src_channel;                                                                        // id_router_029:src_channel -> rsp_xbar_demux_029:sink_channel
	wire          id_router_029_src_ready;                                                                          // rsp_xbar_demux_029:sink_ready -> id_router_029:src_ready
	wire          cmd_xbar_demux_001_src30_ready;                                                                   // CH0_YN3_U_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src30_ready
	wire          id_router_030_src_endofpacket;                                                                    // id_router_030:src_endofpacket -> rsp_xbar_demux_030:sink_endofpacket
	wire          id_router_030_src_valid;                                                                          // id_router_030:src_valid -> rsp_xbar_demux_030:sink_valid
	wire          id_router_030_src_startofpacket;                                                                  // id_router_030:src_startofpacket -> rsp_xbar_demux_030:sink_startofpacket
	wire  [102:0] id_router_030_src_data;                                                                           // id_router_030:src_data -> rsp_xbar_demux_030:sink_data
	wire   [98:0] id_router_030_src_channel;                                                                        // id_router_030:src_channel -> rsp_xbar_demux_030:sink_channel
	wire          id_router_030_src_ready;                                                                          // rsp_xbar_demux_030:sink_ready -> id_router_030:src_ready
	wire          cmd_xbar_demux_001_src31_ready;                                                                   // CH1_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src31_ready
	wire          id_router_031_src_endofpacket;                                                                    // id_router_031:src_endofpacket -> rsp_xbar_demux_031:sink_endofpacket
	wire          id_router_031_src_valid;                                                                          // id_router_031:src_valid -> rsp_xbar_demux_031:sink_valid
	wire          id_router_031_src_startofpacket;                                                                  // id_router_031:src_startofpacket -> rsp_xbar_demux_031:sink_startofpacket
	wire  [102:0] id_router_031_src_data;                                                                           // id_router_031:src_data -> rsp_xbar_demux_031:sink_data
	wire   [98:0] id_router_031_src_channel;                                                                        // id_router_031:src_channel -> rsp_xbar_demux_031:sink_channel
	wire          id_router_031_src_ready;                                                                          // rsp_xbar_demux_031:sink_ready -> id_router_031:src_ready
	wire          cmd_xbar_demux_001_src32_ready;                                                                   // CH1_THRESH_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src32_ready
	wire          id_router_032_src_endofpacket;                                                                    // id_router_032:src_endofpacket -> rsp_xbar_demux_032:sink_endofpacket
	wire          id_router_032_src_valid;                                                                          // id_router_032:src_valid -> rsp_xbar_demux_032:sink_valid
	wire          id_router_032_src_startofpacket;                                                                  // id_router_032:src_startofpacket -> rsp_xbar_demux_032:sink_startofpacket
	wire  [102:0] id_router_032_src_data;                                                                           // id_router_032:src_data -> rsp_xbar_demux_032:sink_data
	wire   [98:0] id_router_032_src_channel;                                                                        // id_router_032:src_channel -> rsp_xbar_demux_032:sink_channel
	wire          id_router_032_src_ready;                                                                          // rsp_xbar_demux_032:sink_ready -> id_router_032:src_ready
	wire          cmd_xbar_demux_001_src33_ready;                                                                   // CH1_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src33_ready
	wire          id_router_033_src_endofpacket;                                                                    // id_router_033:src_endofpacket -> rsp_xbar_demux_033:sink_endofpacket
	wire          id_router_033_src_valid;                                                                          // id_router_033:src_valid -> rsp_xbar_demux_033:sink_valid
	wire          id_router_033_src_startofpacket;                                                                  // id_router_033:src_startofpacket -> rsp_xbar_demux_033:sink_startofpacket
	wire  [102:0] id_router_033_src_data;                                                                           // id_router_033:src_data -> rsp_xbar_demux_033:sink_data
	wire   [98:0] id_router_033_src_channel;                                                                        // id_router_033:src_channel -> rsp_xbar_demux_033:sink_channel
	wire          id_router_033_src_ready;                                                                          // rsp_xbar_demux_033:sink_ready -> id_router_033:src_ready
	wire          cmd_xbar_demux_001_src34_ready;                                                                   // CH1_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src34_ready
	wire          id_router_034_src_endofpacket;                                                                    // id_router_034:src_endofpacket -> rsp_xbar_demux_034:sink_endofpacket
	wire          id_router_034_src_valid;                                                                          // id_router_034:src_valid -> rsp_xbar_demux_034:sink_valid
	wire          id_router_034_src_startofpacket;                                                                  // id_router_034:src_startofpacket -> rsp_xbar_demux_034:sink_startofpacket
	wire  [102:0] id_router_034_src_data;                                                                           // id_router_034:src_data -> rsp_xbar_demux_034:sink_data
	wire   [98:0] id_router_034_src_channel;                                                                        // id_router_034:src_channel -> rsp_xbar_demux_034:sink_channel
	wire          id_router_034_src_ready;                                                                          // rsp_xbar_demux_034:sink_ready -> id_router_034:src_ready
	wire          cmd_xbar_demux_001_src35_ready;                                                                   // CH1_TIME_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src35_ready
	wire          id_router_035_src_endofpacket;                                                                    // id_router_035:src_endofpacket -> rsp_xbar_demux_035:sink_endofpacket
	wire          id_router_035_src_valid;                                                                          // id_router_035:src_valid -> rsp_xbar_demux_035:sink_valid
	wire          id_router_035_src_startofpacket;                                                                  // id_router_035:src_startofpacket -> rsp_xbar_demux_035:sink_startofpacket
	wire  [102:0] id_router_035_src_data;                                                                           // id_router_035:src_data -> rsp_xbar_demux_035:sink_data
	wire   [98:0] id_router_035_src_channel;                                                                        // id_router_035:src_channel -> rsp_xbar_demux_035:sink_channel
	wire          id_router_035_src_ready;                                                                          // rsp_xbar_demux_035:sink_ready -> id_router_035:src_ready
	wire          cmd_xbar_demux_001_src36_ready;                                                                   // CH1_YN1_U_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src36_ready
	wire          id_router_036_src_endofpacket;                                                                    // id_router_036:src_endofpacket -> rsp_xbar_demux_036:sink_endofpacket
	wire          id_router_036_src_valid;                                                                          // id_router_036:src_valid -> rsp_xbar_demux_036:sink_valid
	wire          id_router_036_src_startofpacket;                                                                  // id_router_036:src_startofpacket -> rsp_xbar_demux_036:sink_startofpacket
	wire  [102:0] id_router_036_src_data;                                                                           // id_router_036:src_data -> rsp_xbar_demux_036:sink_data
	wire   [98:0] id_router_036_src_channel;                                                                        // id_router_036:src_channel -> rsp_xbar_demux_036:sink_channel
	wire          id_router_036_src_ready;                                                                          // rsp_xbar_demux_036:sink_ready -> id_router_036:src_ready
	wire          cmd_xbar_demux_001_src37_ready;                                                                   // CH1_YN1_MU_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src37_ready
	wire          id_router_037_src_endofpacket;                                                                    // id_router_037:src_endofpacket -> rsp_xbar_demux_037:sink_endofpacket
	wire          id_router_037_src_valid;                                                                          // id_router_037:src_valid -> rsp_xbar_demux_037:sink_valid
	wire          id_router_037_src_startofpacket;                                                                  // id_router_037:src_startofpacket -> rsp_xbar_demux_037:sink_startofpacket
	wire  [102:0] id_router_037_src_data;                                                                           // id_router_037:src_data -> rsp_xbar_demux_037:sink_data
	wire   [98:0] id_router_037_src_channel;                                                                        // id_router_037:src_channel -> rsp_xbar_demux_037:sink_channel
	wire          id_router_037_src_ready;                                                                          // rsp_xbar_demux_037:sink_ready -> id_router_037:src_ready
	wire          cmd_xbar_demux_001_src38_ready;                                                                   // CH1_YN1_ML_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src38_ready
	wire          id_router_038_src_endofpacket;                                                                    // id_router_038:src_endofpacket -> rsp_xbar_demux_038:sink_endofpacket
	wire          id_router_038_src_valid;                                                                          // id_router_038:src_valid -> rsp_xbar_demux_038:sink_valid
	wire          id_router_038_src_startofpacket;                                                                  // id_router_038:src_startofpacket -> rsp_xbar_demux_038:sink_startofpacket
	wire  [102:0] id_router_038_src_data;                                                                           // id_router_038:src_data -> rsp_xbar_demux_038:sink_data
	wire   [98:0] id_router_038_src_channel;                                                                        // id_router_038:src_channel -> rsp_xbar_demux_038:sink_channel
	wire          id_router_038_src_ready;                                                                          // rsp_xbar_demux_038:sink_ready -> id_router_038:src_ready
	wire          cmd_xbar_demux_001_src39_ready;                                                                   // CH1_YN1_L_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src39_ready
	wire          id_router_039_src_endofpacket;                                                                    // id_router_039:src_endofpacket -> rsp_xbar_demux_039:sink_endofpacket
	wire          id_router_039_src_valid;                                                                          // id_router_039:src_valid -> rsp_xbar_demux_039:sink_valid
	wire          id_router_039_src_startofpacket;                                                                  // id_router_039:src_startofpacket -> rsp_xbar_demux_039:sink_startofpacket
	wire  [102:0] id_router_039_src_data;                                                                           // id_router_039:src_data -> rsp_xbar_demux_039:sink_data
	wire   [98:0] id_router_039_src_channel;                                                                        // id_router_039:src_channel -> rsp_xbar_demux_039:sink_channel
	wire          id_router_039_src_ready;                                                                          // rsp_xbar_demux_039:sink_ready -> id_router_039:src_ready
	wire          cmd_xbar_demux_001_src40_ready;                                                                   // CH1_YN2_U_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src40_ready
	wire          id_router_040_src_endofpacket;                                                                    // id_router_040:src_endofpacket -> rsp_xbar_demux_040:sink_endofpacket
	wire          id_router_040_src_valid;                                                                          // id_router_040:src_valid -> rsp_xbar_demux_040:sink_valid
	wire          id_router_040_src_startofpacket;                                                                  // id_router_040:src_startofpacket -> rsp_xbar_demux_040:sink_startofpacket
	wire  [102:0] id_router_040_src_data;                                                                           // id_router_040:src_data -> rsp_xbar_demux_040:sink_data
	wire   [98:0] id_router_040_src_channel;                                                                        // id_router_040:src_channel -> rsp_xbar_demux_040:sink_channel
	wire          id_router_040_src_ready;                                                                          // rsp_xbar_demux_040:sink_ready -> id_router_040:src_ready
	wire          cmd_xbar_demux_001_src41_ready;                                                                   // CH1_YN2_MU_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src41_ready
	wire          id_router_041_src_endofpacket;                                                                    // id_router_041:src_endofpacket -> rsp_xbar_demux_041:sink_endofpacket
	wire          id_router_041_src_valid;                                                                          // id_router_041:src_valid -> rsp_xbar_demux_041:sink_valid
	wire          id_router_041_src_startofpacket;                                                                  // id_router_041:src_startofpacket -> rsp_xbar_demux_041:sink_startofpacket
	wire  [102:0] id_router_041_src_data;                                                                           // id_router_041:src_data -> rsp_xbar_demux_041:sink_data
	wire   [98:0] id_router_041_src_channel;                                                                        // id_router_041:src_channel -> rsp_xbar_demux_041:sink_channel
	wire          id_router_041_src_ready;                                                                          // rsp_xbar_demux_041:sink_ready -> id_router_041:src_ready
	wire          cmd_xbar_demux_001_src42_ready;                                                                   // CH1_YN2_ML_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src42_ready
	wire          id_router_042_src_endofpacket;                                                                    // id_router_042:src_endofpacket -> rsp_xbar_demux_042:sink_endofpacket
	wire          id_router_042_src_valid;                                                                          // id_router_042:src_valid -> rsp_xbar_demux_042:sink_valid
	wire          id_router_042_src_startofpacket;                                                                  // id_router_042:src_startofpacket -> rsp_xbar_demux_042:sink_startofpacket
	wire  [102:0] id_router_042_src_data;                                                                           // id_router_042:src_data -> rsp_xbar_demux_042:sink_data
	wire   [98:0] id_router_042_src_channel;                                                                        // id_router_042:src_channel -> rsp_xbar_demux_042:sink_channel
	wire          id_router_042_src_ready;                                                                          // rsp_xbar_demux_042:sink_ready -> id_router_042:src_ready
	wire          cmd_xbar_demux_001_src43_ready;                                                                   // CH1_YN2_L_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src43_ready
	wire          id_router_043_src_endofpacket;                                                                    // id_router_043:src_endofpacket -> rsp_xbar_demux_043:sink_endofpacket
	wire          id_router_043_src_valid;                                                                          // id_router_043:src_valid -> rsp_xbar_demux_043:sink_valid
	wire          id_router_043_src_startofpacket;                                                                  // id_router_043:src_startofpacket -> rsp_xbar_demux_043:sink_startofpacket
	wire  [102:0] id_router_043_src_data;                                                                           // id_router_043:src_data -> rsp_xbar_demux_043:sink_data
	wire   [98:0] id_router_043_src_channel;                                                                        // id_router_043:src_channel -> rsp_xbar_demux_043:sink_channel
	wire          id_router_043_src_ready;                                                                          // rsp_xbar_demux_043:sink_ready -> id_router_043:src_ready
	wire          cmd_xbar_demux_001_src44_ready;                                                                   // CH1_YN3_U_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src44_ready
	wire          id_router_044_src_endofpacket;                                                                    // id_router_044:src_endofpacket -> rsp_xbar_demux_044:sink_endofpacket
	wire          id_router_044_src_valid;                                                                          // id_router_044:src_valid -> rsp_xbar_demux_044:sink_valid
	wire          id_router_044_src_startofpacket;                                                                  // id_router_044:src_startofpacket -> rsp_xbar_demux_044:sink_startofpacket
	wire  [102:0] id_router_044_src_data;                                                                           // id_router_044:src_data -> rsp_xbar_demux_044:sink_data
	wire   [98:0] id_router_044_src_channel;                                                                        // id_router_044:src_channel -> rsp_xbar_demux_044:sink_channel
	wire          id_router_044_src_ready;                                                                          // rsp_xbar_demux_044:sink_ready -> id_router_044:src_ready
	wire          cmd_xbar_demux_001_src45_ready;                                                                   // CH1_YN3_MU_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src45_ready
	wire          id_router_045_src_endofpacket;                                                                    // id_router_045:src_endofpacket -> rsp_xbar_demux_045:sink_endofpacket
	wire          id_router_045_src_valid;                                                                          // id_router_045:src_valid -> rsp_xbar_demux_045:sink_valid
	wire          id_router_045_src_startofpacket;                                                                  // id_router_045:src_startofpacket -> rsp_xbar_demux_045:sink_startofpacket
	wire  [102:0] id_router_045_src_data;                                                                           // id_router_045:src_data -> rsp_xbar_demux_045:sink_data
	wire   [98:0] id_router_045_src_channel;                                                                        // id_router_045:src_channel -> rsp_xbar_demux_045:sink_channel
	wire          id_router_045_src_ready;                                                                          // rsp_xbar_demux_045:sink_ready -> id_router_045:src_ready
	wire          cmd_xbar_demux_001_src46_ready;                                                                   // CH1_YN3_ML_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src46_ready
	wire          id_router_046_src_endofpacket;                                                                    // id_router_046:src_endofpacket -> rsp_xbar_demux_046:sink_endofpacket
	wire          id_router_046_src_valid;                                                                          // id_router_046:src_valid -> rsp_xbar_demux_046:sink_valid
	wire          id_router_046_src_startofpacket;                                                                  // id_router_046:src_startofpacket -> rsp_xbar_demux_046:sink_startofpacket
	wire  [102:0] id_router_046_src_data;                                                                           // id_router_046:src_data -> rsp_xbar_demux_046:sink_data
	wire   [98:0] id_router_046_src_channel;                                                                        // id_router_046:src_channel -> rsp_xbar_demux_046:sink_channel
	wire          id_router_046_src_ready;                                                                          // rsp_xbar_demux_046:sink_ready -> id_router_046:src_ready
	wire          cmd_xbar_demux_001_src47_ready;                                                                   // CH1_YN3_L_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src47_ready
	wire          id_router_047_src_endofpacket;                                                                    // id_router_047:src_endofpacket -> rsp_xbar_demux_047:sink_endofpacket
	wire          id_router_047_src_valid;                                                                          // id_router_047:src_valid -> rsp_xbar_demux_047:sink_valid
	wire          id_router_047_src_startofpacket;                                                                  // id_router_047:src_startofpacket -> rsp_xbar_demux_047:sink_startofpacket
	wire  [102:0] id_router_047_src_data;                                                                           // id_router_047:src_data -> rsp_xbar_demux_047:sink_data
	wire   [98:0] id_router_047_src_channel;                                                                        // id_router_047:src_channel -> rsp_xbar_demux_047:sink_channel
	wire          id_router_047_src_ready;                                                                          // rsp_xbar_demux_047:sink_ready -> id_router_047:src_ready
	wire          cmd_xbar_demux_001_src48_ready;                                                                   // CH2_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src48_ready
	wire          id_router_048_src_endofpacket;                                                                    // id_router_048:src_endofpacket -> rsp_xbar_demux_048:sink_endofpacket
	wire          id_router_048_src_valid;                                                                          // id_router_048:src_valid -> rsp_xbar_demux_048:sink_valid
	wire          id_router_048_src_startofpacket;                                                                  // id_router_048:src_startofpacket -> rsp_xbar_demux_048:sink_startofpacket
	wire  [102:0] id_router_048_src_data;                                                                           // id_router_048:src_data -> rsp_xbar_demux_048:sink_data
	wire   [98:0] id_router_048_src_channel;                                                                        // id_router_048:src_channel -> rsp_xbar_demux_048:sink_channel
	wire          id_router_048_src_ready;                                                                          // rsp_xbar_demux_048:sink_ready -> id_router_048:src_ready
	wire          cmd_xbar_demux_001_src49_ready;                                                                   // CH2_THRESH_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src49_ready
	wire          id_router_049_src_endofpacket;                                                                    // id_router_049:src_endofpacket -> rsp_xbar_demux_049:sink_endofpacket
	wire          id_router_049_src_valid;                                                                          // id_router_049:src_valid -> rsp_xbar_demux_049:sink_valid
	wire          id_router_049_src_startofpacket;                                                                  // id_router_049:src_startofpacket -> rsp_xbar_demux_049:sink_startofpacket
	wire  [102:0] id_router_049_src_data;                                                                           // id_router_049:src_data -> rsp_xbar_demux_049:sink_data
	wire   [98:0] id_router_049_src_channel;                                                                        // id_router_049:src_channel -> rsp_xbar_demux_049:sink_channel
	wire          id_router_049_src_ready;                                                                          // rsp_xbar_demux_049:sink_ready -> id_router_049:src_ready
	wire          cmd_xbar_demux_001_src50_ready;                                                                   // CH2_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src50_ready
	wire          id_router_050_src_endofpacket;                                                                    // id_router_050:src_endofpacket -> rsp_xbar_demux_050:sink_endofpacket
	wire          id_router_050_src_valid;                                                                          // id_router_050:src_valid -> rsp_xbar_demux_050:sink_valid
	wire          id_router_050_src_startofpacket;                                                                  // id_router_050:src_startofpacket -> rsp_xbar_demux_050:sink_startofpacket
	wire  [102:0] id_router_050_src_data;                                                                           // id_router_050:src_data -> rsp_xbar_demux_050:sink_data
	wire   [98:0] id_router_050_src_channel;                                                                        // id_router_050:src_channel -> rsp_xbar_demux_050:sink_channel
	wire          id_router_050_src_ready;                                                                          // rsp_xbar_demux_050:sink_ready -> id_router_050:src_ready
	wire          cmd_xbar_demux_001_src51_ready;                                                                   // CH2_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src51_ready
	wire          id_router_051_src_endofpacket;                                                                    // id_router_051:src_endofpacket -> rsp_xbar_demux_051:sink_endofpacket
	wire          id_router_051_src_valid;                                                                          // id_router_051:src_valid -> rsp_xbar_demux_051:sink_valid
	wire          id_router_051_src_startofpacket;                                                                  // id_router_051:src_startofpacket -> rsp_xbar_demux_051:sink_startofpacket
	wire  [102:0] id_router_051_src_data;                                                                           // id_router_051:src_data -> rsp_xbar_demux_051:sink_data
	wire   [98:0] id_router_051_src_channel;                                                                        // id_router_051:src_channel -> rsp_xbar_demux_051:sink_channel
	wire          id_router_051_src_ready;                                                                          // rsp_xbar_demux_051:sink_ready -> id_router_051:src_ready
	wire          cmd_xbar_demux_001_src52_ready;                                                                   // CH2_TIME_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src52_ready
	wire          id_router_052_src_endofpacket;                                                                    // id_router_052:src_endofpacket -> rsp_xbar_demux_052:sink_endofpacket
	wire          id_router_052_src_valid;                                                                          // id_router_052:src_valid -> rsp_xbar_demux_052:sink_valid
	wire          id_router_052_src_startofpacket;                                                                  // id_router_052:src_startofpacket -> rsp_xbar_demux_052:sink_startofpacket
	wire  [102:0] id_router_052_src_data;                                                                           // id_router_052:src_data -> rsp_xbar_demux_052:sink_data
	wire   [98:0] id_router_052_src_channel;                                                                        // id_router_052:src_channel -> rsp_xbar_demux_052:sink_channel
	wire          id_router_052_src_ready;                                                                          // rsp_xbar_demux_052:sink_ready -> id_router_052:src_ready
	wire          cmd_xbar_demux_001_src53_ready;                                                                   // CH2_YN1_U_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src53_ready
	wire          id_router_053_src_endofpacket;                                                                    // id_router_053:src_endofpacket -> rsp_xbar_demux_053:sink_endofpacket
	wire          id_router_053_src_valid;                                                                          // id_router_053:src_valid -> rsp_xbar_demux_053:sink_valid
	wire          id_router_053_src_startofpacket;                                                                  // id_router_053:src_startofpacket -> rsp_xbar_demux_053:sink_startofpacket
	wire  [102:0] id_router_053_src_data;                                                                           // id_router_053:src_data -> rsp_xbar_demux_053:sink_data
	wire   [98:0] id_router_053_src_channel;                                                                        // id_router_053:src_channel -> rsp_xbar_demux_053:sink_channel
	wire          id_router_053_src_ready;                                                                          // rsp_xbar_demux_053:sink_ready -> id_router_053:src_ready
	wire          cmd_xbar_demux_001_src54_ready;                                                                   // CH2_YN1_MU_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src54_ready
	wire          id_router_054_src_endofpacket;                                                                    // id_router_054:src_endofpacket -> rsp_xbar_demux_054:sink_endofpacket
	wire          id_router_054_src_valid;                                                                          // id_router_054:src_valid -> rsp_xbar_demux_054:sink_valid
	wire          id_router_054_src_startofpacket;                                                                  // id_router_054:src_startofpacket -> rsp_xbar_demux_054:sink_startofpacket
	wire  [102:0] id_router_054_src_data;                                                                           // id_router_054:src_data -> rsp_xbar_demux_054:sink_data
	wire   [98:0] id_router_054_src_channel;                                                                        // id_router_054:src_channel -> rsp_xbar_demux_054:sink_channel
	wire          id_router_054_src_ready;                                                                          // rsp_xbar_demux_054:sink_ready -> id_router_054:src_ready
	wire          cmd_xbar_demux_001_src55_ready;                                                                   // CH2_YN1_ML_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src55_ready
	wire          id_router_055_src_endofpacket;                                                                    // id_router_055:src_endofpacket -> rsp_xbar_demux_055:sink_endofpacket
	wire          id_router_055_src_valid;                                                                          // id_router_055:src_valid -> rsp_xbar_demux_055:sink_valid
	wire          id_router_055_src_startofpacket;                                                                  // id_router_055:src_startofpacket -> rsp_xbar_demux_055:sink_startofpacket
	wire  [102:0] id_router_055_src_data;                                                                           // id_router_055:src_data -> rsp_xbar_demux_055:sink_data
	wire   [98:0] id_router_055_src_channel;                                                                        // id_router_055:src_channel -> rsp_xbar_demux_055:sink_channel
	wire          id_router_055_src_ready;                                                                          // rsp_xbar_demux_055:sink_ready -> id_router_055:src_ready
	wire          cmd_xbar_demux_001_src56_ready;                                                                   // CH2_YN1_L_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src56_ready
	wire          id_router_056_src_endofpacket;                                                                    // id_router_056:src_endofpacket -> rsp_xbar_demux_056:sink_endofpacket
	wire          id_router_056_src_valid;                                                                          // id_router_056:src_valid -> rsp_xbar_demux_056:sink_valid
	wire          id_router_056_src_startofpacket;                                                                  // id_router_056:src_startofpacket -> rsp_xbar_demux_056:sink_startofpacket
	wire  [102:0] id_router_056_src_data;                                                                           // id_router_056:src_data -> rsp_xbar_demux_056:sink_data
	wire   [98:0] id_router_056_src_channel;                                                                        // id_router_056:src_channel -> rsp_xbar_demux_056:sink_channel
	wire          id_router_056_src_ready;                                                                          // rsp_xbar_demux_056:sink_ready -> id_router_056:src_ready
	wire          cmd_xbar_demux_001_src57_ready;                                                                   // CH2_YN2_U_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src57_ready
	wire          id_router_057_src_endofpacket;                                                                    // id_router_057:src_endofpacket -> rsp_xbar_demux_057:sink_endofpacket
	wire          id_router_057_src_valid;                                                                          // id_router_057:src_valid -> rsp_xbar_demux_057:sink_valid
	wire          id_router_057_src_startofpacket;                                                                  // id_router_057:src_startofpacket -> rsp_xbar_demux_057:sink_startofpacket
	wire  [102:0] id_router_057_src_data;                                                                           // id_router_057:src_data -> rsp_xbar_demux_057:sink_data
	wire   [98:0] id_router_057_src_channel;                                                                        // id_router_057:src_channel -> rsp_xbar_demux_057:sink_channel
	wire          id_router_057_src_ready;                                                                          // rsp_xbar_demux_057:sink_ready -> id_router_057:src_ready
	wire          cmd_xbar_demux_001_src58_ready;                                                                   // CH2_YN2_MU_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src58_ready
	wire          id_router_058_src_endofpacket;                                                                    // id_router_058:src_endofpacket -> rsp_xbar_demux_058:sink_endofpacket
	wire          id_router_058_src_valid;                                                                          // id_router_058:src_valid -> rsp_xbar_demux_058:sink_valid
	wire          id_router_058_src_startofpacket;                                                                  // id_router_058:src_startofpacket -> rsp_xbar_demux_058:sink_startofpacket
	wire  [102:0] id_router_058_src_data;                                                                           // id_router_058:src_data -> rsp_xbar_demux_058:sink_data
	wire   [98:0] id_router_058_src_channel;                                                                        // id_router_058:src_channel -> rsp_xbar_demux_058:sink_channel
	wire          id_router_058_src_ready;                                                                          // rsp_xbar_demux_058:sink_ready -> id_router_058:src_ready
	wire          cmd_xbar_demux_001_src59_ready;                                                                   // CH2_YN2_ML_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src59_ready
	wire          id_router_059_src_endofpacket;                                                                    // id_router_059:src_endofpacket -> rsp_xbar_demux_059:sink_endofpacket
	wire          id_router_059_src_valid;                                                                          // id_router_059:src_valid -> rsp_xbar_demux_059:sink_valid
	wire          id_router_059_src_startofpacket;                                                                  // id_router_059:src_startofpacket -> rsp_xbar_demux_059:sink_startofpacket
	wire  [102:0] id_router_059_src_data;                                                                           // id_router_059:src_data -> rsp_xbar_demux_059:sink_data
	wire   [98:0] id_router_059_src_channel;                                                                        // id_router_059:src_channel -> rsp_xbar_demux_059:sink_channel
	wire          id_router_059_src_ready;                                                                          // rsp_xbar_demux_059:sink_ready -> id_router_059:src_ready
	wire          cmd_xbar_demux_001_src60_ready;                                                                   // CH2_YN2_L_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src60_ready
	wire          id_router_060_src_endofpacket;                                                                    // id_router_060:src_endofpacket -> rsp_xbar_demux_060:sink_endofpacket
	wire          id_router_060_src_valid;                                                                          // id_router_060:src_valid -> rsp_xbar_demux_060:sink_valid
	wire          id_router_060_src_startofpacket;                                                                  // id_router_060:src_startofpacket -> rsp_xbar_demux_060:sink_startofpacket
	wire  [102:0] id_router_060_src_data;                                                                           // id_router_060:src_data -> rsp_xbar_demux_060:sink_data
	wire   [98:0] id_router_060_src_channel;                                                                        // id_router_060:src_channel -> rsp_xbar_demux_060:sink_channel
	wire          id_router_060_src_ready;                                                                          // rsp_xbar_demux_060:sink_ready -> id_router_060:src_ready
	wire          cmd_xbar_demux_001_src61_ready;                                                                   // CH2_YN3_U_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src61_ready
	wire          id_router_061_src_endofpacket;                                                                    // id_router_061:src_endofpacket -> rsp_xbar_demux_061:sink_endofpacket
	wire          id_router_061_src_valid;                                                                          // id_router_061:src_valid -> rsp_xbar_demux_061:sink_valid
	wire          id_router_061_src_startofpacket;                                                                  // id_router_061:src_startofpacket -> rsp_xbar_demux_061:sink_startofpacket
	wire  [102:0] id_router_061_src_data;                                                                           // id_router_061:src_data -> rsp_xbar_demux_061:sink_data
	wire   [98:0] id_router_061_src_channel;                                                                        // id_router_061:src_channel -> rsp_xbar_demux_061:sink_channel
	wire          id_router_061_src_ready;                                                                          // rsp_xbar_demux_061:sink_ready -> id_router_061:src_ready
	wire          cmd_xbar_demux_001_src62_ready;                                                                   // CH2_YN3_MU_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src62_ready
	wire          id_router_062_src_endofpacket;                                                                    // id_router_062:src_endofpacket -> rsp_xbar_demux_062:sink_endofpacket
	wire          id_router_062_src_valid;                                                                          // id_router_062:src_valid -> rsp_xbar_demux_062:sink_valid
	wire          id_router_062_src_startofpacket;                                                                  // id_router_062:src_startofpacket -> rsp_xbar_demux_062:sink_startofpacket
	wire  [102:0] id_router_062_src_data;                                                                           // id_router_062:src_data -> rsp_xbar_demux_062:sink_data
	wire   [98:0] id_router_062_src_channel;                                                                        // id_router_062:src_channel -> rsp_xbar_demux_062:sink_channel
	wire          id_router_062_src_ready;                                                                          // rsp_xbar_demux_062:sink_ready -> id_router_062:src_ready
	wire          cmd_xbar_demux_001_src63_ready;                                                                   // CH2_YN3_ML_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src63_ready
	wire          id_router_063_src_endofpacket;                                                                    // id_router_063:src_endofpacket -> rsp_xbar_demux_063:sink_endofpacket
	wire          id_router_063_src_valid;                                                                          // id_router_063:src_valid -> rsp_xbar_demux_063:sink_valid
	wire          id_router_063_src_startofpacket;                                                                  // id_router_063:src_startofpacket -> rsp_xbar_demux_063:sink_startofpacket
	wire  [102:0] id_router_063_src_data;                                                                           // id_router_063:src_data -> rsp_xbar_demux_063:sink_data
	wire   [98:0] id_router_063_src_channel;                                                                        // id_router_063:src_channel -> rsp_xbar_demux_063:sink_channel
	wire          id_router_063_src_ready;                                                                          // rsp_xbar_demux_063:sink_ready -> id_router_063:src_ready
	wire          cmd_xbar_demux_001_src64_ready;                                                                   // CH2_YN3_L_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src64_ready
	wire          id_router_064_src_endofpacket;                                                                    // id_router_064:src_endofpacket -> rsp_xbar_demux_064:sink_endofpacket
	wire          id_router_064_src_valid;                                                                          // id_router_064:src_valid -> rsp_xbar_demux_064:sink_valid
	wire          id_router_064_src_startofpacket;                                                                  // id_router_064:src_startofpacket -> rsp_xbar_demux_064:sink_startofpacket
	wire  [102:0] id_router_064_src_data;                                                                           // id_router_064:src_data -> rsp_xbar_demux_064:sink_data
	wire   [98:0] id_router_064_src_channel;                                                                        // id_router_064:src_channel -> rsp_xbar_demux_064:sink_channel
	wire          id_router_064_src_ready;                                                                          // rsp_xbar_demux_064:sink_ready -> id_router_064:src_ready
	wire          cmd_xbar_demux_001_src65_ready;                                                                   // CH3_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src65_ready
	wire          id_router_065_src_endofpacket;                                                                    // id_router_065:src_endofpacket -> rsp_xbar_demux_065:sink_endofpacket
	wire          id_router_065_src_valid;                                                                          // id_router_065:src_valid -> rsp_xbar_demux_065:sink_valid
	wire          id_router_065_src_startofpacket;                                                                  // id_router_065:src_startofpacket -> rsp_xbar_demux_065:sink_startofpacket
	wire  [102:0] id_router_065_src_data;                                                                           // id_router_065:src_data -> rsp_xbar_demux_065:sink_data
	wire   [98:0] id_router_065_src_channel;                                                                        // id_router_065:src_channel -> rsp_xbar_demux_065:sink_channel
	wire          id_router_065_src_ready;                                                                          // rsp_xbar_demux_065:sink_ready -> id_router_065:src_ready
	wire          cmd_xbar_demux_001_src66_ready;                                                                   // CH3_THRESH_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src66_ready
	wire          id_router_066_src_endofpacket;                                                                    // id_router_066:src_endofpacket -> rsp_xbar_demux_066:sink_endofpacket
	wire          id_router_066_src_valid;                                                                          // id_router_066:src_valid -> rsp_xbar_demux_066:sink_valid
	wire          id_router_066_src_startofpacket;                                                                  // id_router_066:src_startofpacket -> rsp_xbar_demux_066:sink_startofpacket
	wire  [102:0] id_router_066_src_data;                                                                           // id_router_066:src_data -> rsp_xbar_demux_066:sink_data
	wire   [98:0] id_router_066_src_channel;                                                                        // id_router_066:src_channel -> rsp_xbar_demux_066:sink_channel
	wire          id_router_066_src_ready;                                                                          // rsp_xbar_demux_066:sink_ready -> id_router_066:src_ready
	wire          cmd_xbar_demux_001_src67_ready;                                                                   // CH3_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src67_ready
	wire          id_router_067_src_endofpacket;                                                                    // id_router_067:src_endofpacket -> rsp_xbar_demux_067:sink_endofpacket
	wire          id_router_067_src_valid;                                                                          // id_router_067:src_valid -> rsp_xbar_demux_067:sink_valid
	wire          id_router_067_src_startofpacket;                                                                  // id_router_067:src_startofpacket -> rsp_xbar_demux_067:sink_startofpacket
	wire  [102:0] id_router_067_src_data;                                                                           // id_router_067:src_data -> rsp_xbar_demux_067:sink_data
	wire   [98:0] id_router_067_src_channel;                                                                        // id_router_067:src_channel -> rsp_xbar_demux_067:sink_channel
	wire          id_router_067_src_ready;                                                                          // rsp_xbar_demux_067:sink_ready -> id_router_067:src_ready
	wire          cmd_xbar_demux_001_src68_ready;                                                                   // CH3_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src68_ready
	wire          id_router_068_src_endofpacket;                                                                    // id_router_068:src_endofpacket -> rsp_xbar_demux_068:sink_endofpacket
	wire          id_router_068_src_valid;                                                                          // id_router_068:src_valid -> rsp_xbar_demux_068:sink_valid
	wire          id_router_068_src_startofpacket;                                                                  // id_router_068:src_startofpacket -> rsp_xbar_demux_068:sink_startofpacket
	wire  [102:0] id_router_068_src_data;                                                                           // id_router_068:src_data -> rsp_xbar_demux_068:sink_data
	wire   [98:0] id_router_068_src_channel;                                                                        // id_router_068:src_channel -> rsp_xbar_demux_068:sink_channel
	wire          id_router_068_src_ready;                                                                          // rsp_xbar_demux_068:sink_ready -> id_router_068:src_ready
	wire          cmd_xbar_demux_001_src69_ready;                                                                   // CH3_YN1_U_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src69_ready
	wire          id_router_069_src_endofpacket;                                                                    // id_router_069:src_endofpacket -> rsp_xbar_demux_069:sink_endofpacket
	wire          id_router_069_src_valid;                                                                          // id_router_069:src_valid -> rsp_xbar_demux_069:sink_valid
	wire          id_router_069_src_startofpacket;                                                                  // id_router_069:src_startofpacket -> rsp_xbar_demux_069:sink_startofpacket
	wire  [102:0] id_router_069_src_data;                                                                           // id_router_069:src_data -> rsp_xbar_demux_069:sink_data
	wire   [98:0] id_router_069_src_channel;                                                                        // id_router_069:src_channel -> rsp_xbar_demux_069:sink_channel
	wire          id_router_069_src_ready;                                                                          // rsp_xbar_demux_069:sink_ready -> id_router_069:src_ready
	wire          cmd_xbar_demux_001_src70_ready;                                                                   // CH3_TIME_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src70_ready
	wire          id_router_070_src_endofpacket;                                                                    // id_router_070:src_endofpacket -> rsp_xbar_demux_070:sink_endofpacket
	wire          id_router_070_src_valid;                                                                          // id_router_070:src_valid -> rsp_xbar_demux_070:sink_valid
	wire          id_router_070_src_startofpacket;                                                                  // id_router_070:src_startofpacket -> rsp_xbar_demux_070:sink_startofpacket
	wire  [102:0] id_router_070_src_data;                                                                           // id_router_070:src_data -> rsp_xbar_demux_070:sink_data
	wire   [98:0] id_router_070_src_channel;                                                                        // id_router_070:src_channel -> rsp_xbar_demux_070:sink_channel
	wire          id_router_070_src_ready;                                                                          // rsp_xbar_demux_070:sink_ready -> id_router_070:src_ready
	wire          cmd_xbar_demux_001_src71_ready;                                                                   // CH3_YN3_L_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src71_ready
	wire          id_router_071_src_endofpacket;                                                                    // id_router_071:src_endofpacket -> rsp_xbar_demux_071:sink_endofpacket
	wire          id_router_071_src_valid;                                                                          // id_router_071:src_valid -> rsp_xbar_demux_071:sink_valid
	wire          id_router_071_src_startofpacket;                                                                  // id_router_071:src_startofpacket -> rsp_xbar_demux_071:sink_startofpacket
	wire  [102:0] id_router_071_src_data;                                                                           // id_router_071:src_data -> rsp_xbar_demux_071:sink_data
	wire   [98:0] id_router_071_src_channel;                                                                        // id_router_071:src_channel -> rsp_xbar_demux_071:sink_channel
	wire          id_router_071_src_ready;                                                                          // rsp_xbar_demux_071:sink_ready -> id_router_071:src_ready
	wire          cmd_xbar_demux_001_src72_ready;                                                                   // CH3_YN3_ML_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src72_ready
	wire          id_router_072_src_endofpacket;                                                                    // id_router_072:src_endofpacket -> rsp_xbar_demux_072:sink_endofpacket
	wire          id_router_072_src_valid;                                                                          // id_router_072:src_valid -> rsp_xbar_demux_072:sink_valid
	wire          id_router_072_src_startofpacket;                                                                  // id_router_072:src_startofpacket -> rsp_xbar_demux_072:sink_startofpacket
	wire  [102:0] id_router_072_src_data;                                                                           // id_router_072:src_data -> rsp_xbar_demux_072:sink_data
	wire   [98:0] id_router_072_src_channel;                                                                        // id_router_072:src_channel -> rsp_xbar_demux_072:sink_channel
	wire          id_router_072_src_ready;                                                                          // rsp_xbar_demux_072:sink_ready -> id_router_072:src_ready
	wire          cmd_xbar_demux_001_src73_ready;                                                                   // CH3_YN3_MU_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src73_ready
	wire          id_router_073_src_endofpacket;                                                                    // id_router_073:src_endofpacket -> rsp_xbar_demux_073:sink_endofpacket
	wire          id_router_073_src_valid;                                                                          // id_router_073:src_valid -> rsp_xbar_demux_073:sink_valid
	wire          id_router_073_src_startofpacket;                                                                  // id_router_073:src_startofpacket -> rsp_xbar_demux_073:sink_startofpacket
	wire  [102:0] id_router_073_src_data;                                                                           // id_router_073:src_data -> rsp_xbar_demux_073:sink_data
	wire   [98:0] id_router_073_src_channel;                                                                        // id_router_073:src_channel -> rsp_xbar_demux_073:sink_channel
	wire          id_router_073_src_ready;                                                                          // rsp_xbar_demux_073:sink_ready -> id_router_073:src_ready
	wire          cmd_xbar_demux_001_src74_ready;                                                                   // CH3_YN3_U_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src74_ready
	wire          id_router_074_src_endofpacket;                                                                    // id_router_074:src_endofpacket -> rsp_xbar_demux_074:sink_endofpacket
	wire          id_router_074_src_valid;                                                                          // id_router_074:src_valid -> rsp_xbar_demux_074:sink_valid
	wire          id_router_074_src_startofpacket;                                                                  // id_router_074:src_startofpacket -> rsp_xbar_demux_074:sink_startofpacket
	wire  [102:0] id_router_074_src_data;                                                                           // id_router_074:src_data -> rsp_xbar_demux_074:sink_data
	wire   [98:0] id_router_074_src_channel;                                                                        // id_router_074:src_channel -> rsp_xbar_demux_074:sink_channel
	wire          id_router_074_src_ready;                                                                          // rsp_xbar_demux_074:sink_ready -> id_router_074:src_ready
	wire          cmd_xbar_demux_001_src75_ready;                                                                   // CH3_YN2_L_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src75_ready
	wire          id_router_075_src_endofpacket;                                                                    // id_router_075:src_endofpacket -> rsp_xbar_demux_075:sink_endofpacket
	wire          id_router_075_src_valid;                                                                          // id_router_075:src_valid -> rsp_xbar_demux_075:sink_valid
	wire          id_router_075_src_startofpacket;                                                                  // id_router_075:src_startofpacket -> rsp_xbar_demux_075:sink_startofpacket
	wire  [102:0] id_router_075_src_data;                                                                           // id_router_075:src_data -> rsp_xbar_demux_075:sink_data
	wire   [98:0] id_router_075_src_channel;                                                                        // id_router_075:src_channel -> rsp_xbar_demux_075:sink_channel
	wire          id_router_075_src_ready;                                                                          // rsp_xbar_demux_075:sink_ready -> id_router_075:src_ready
	wire          cmd_xbar_demux_001_src76_ready;                                                                   // CH3_YN2_ML_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src76_ready
	wire          id_router_076_src_endofpacket;                                                                    // id_router_076:src_endofpacket -> rsp_xbar_demux_076:sink_endofpacket
	wire          id_router_076_src_valid;                                                                          // id_router_076:src_valid -> rsp_xbar_demux_076:sink_valid
	wire          id_router_076_src_startofpacket;                                                                  // id_router_076:src_startofpacket -> rsp_xbar_demux_076:sink_startofpacket
	wire  [102:0] id_router_076_src_data;                                                                           // id_router_076:src_data -> rsp_xbar_demux_076:sink_data
	wire   [98:0] id_router_076_src_channel;                                                                        // id_router_076:src_channel -> rsp_xbar_demux_076:sink_channel
	wire          id_router_076_src_ready;                                                                          // rsp_xbar_demux_076:sink_ready -> id_router_076:src_ready
	wire          cmd_xbar_demux_001_src77_ready;                                                                   // CH3_YN2_MU_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src77_ready
	wire          id_router_077_src_endofpacket;                                                                    // id_router_077:src_endofpacket -> rsp_xbar_demux_077:sink_endofpacket
	wire          id_router_077_src_valid;                                                                          // id_router_077:src_valid -> rsp_xbar_demux_077:sink_valid
	wire          id_router_077_src_startofpacket;                                                                  // id_router_077:src_startofpacket -> rsp_xbar_demux_077:sink_startofpacket
	wire  [102:0] id_router_077_src_data;                                                                           // id_router_077:src_data -> rsp_xbar_demux_077:sink_data
	wire   [98:0] id_router_077_src_channel;                                                                        // id_router_077:src_channel -> rsp_xbar_demux_077:sink_channel
	wire          id_router_077_src_ready;                                                                          // rsp_xbar_demux_077:sink_ready -> id_router_077:src_ready
	wire          cmd_xbar_demux_001_src78_ready;                                                                   // CH3_YN2_U_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src78_ready
	wire          id_router_078_src_endofpacket;                                                                    // id_router_078:src_endofpacket -> rsp_xbar_demux_078:sink_endofpacket
	wire          id_router_078_src_valid;                                                                          // id_router_078:src_valid -> rsp_xbar_demux_078:sink_valid
	wire          id_router_078_src_startofpacket;                                                                  // id_router_078:src_startofpacket -> rsp_xbar_demux_078:sink_startofpacket
	wire  [102:0] id_router_078_src_data;                                                                           // id_router_078:src_data -> rsp_xbar_demux_078:sink_data
	wire   [98:0] id_router_078_src_channel;                                                                        // id_router_078:src_channel -> rsp_xbar_demux_078:sink_channel
	wire          id_router_078_src_ready;                                                                          // rsp_xbar_demux_078:sink_ready -> id_router_078:src_ready
	wire          cmd_xbar_demux_001_src79_ready;                                                                   // CH3_YN1_L_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src79_ready
	wire          id_router_079_src_endofpacket;                                                                    // id_router_079:src_endofpacket -> rsp_xbar_demux_079:sink_endofpacket
	wire          id_router_079_src_valid;                                                                          // id_router_079:src_valid -> rsp_xbar_demux_079:sink_valid
	wire          id_router_079_src_startofpacket;                                                                  // id_router_079:src_startofpacket -> rsp_xbar_demux_079:sink_startofpacket
	wire  [102:0] id_router_079_src_data;                                                                           // id_router_079:src_data -> rsp_xbar_demux_079:sink_data
	wire   [98:0] id_router_079_src_channel;                                                                        // id_router_079:src_channel -> rsp_xbar_demux_079:sink_channel
	wire          id_router_079_src_ready;                                                                          // rsp_xbar_demux_079:sink_ready -> id_router_079:src_ready
	wire          cmd_xbar_demux_001_src80_ready;                                                                   // CH3_YN1_MU_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src80_ready
	wire          id_router_080_src_endofpacket;                                                                    // id_router_080:src_endofpacket -> rsp_xbar_demux_080:sink_endofpacket
	wire          id_router_080_src_valid;                                                                          // id_router_080:src_valid -> rsp_xbar_demux_080:sink_valid
	wire          id_router_080_src_startofpacket;                                                                  // id_router_080:src_startofpacket -> rsp_xbar_demux_080:sink_startofpacket
	wire  [102:0] id_router_080_src_data;                                                                           // id_router_080:src_data -> rsp_xbar_demux_080:sink_data
	wire   [98:0] id_router_080_src_channel;                                                                        // id_router_080:src_channel -> rsp_xbar_demux_080:sink_channel
	wire          id_router_080_src_ready;                                                                          // rsp_xbar_demux_080:sink_ready -> id_router_080:src_ready
	wire          cmd_xbar_demux_001_src81_ready;                                                                   // CH3_YN1_ML_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src81_ready
	wire          id_router_081_src_endofpacket;                                                                    // id_router_081:src_endofpacket -> rsp_xbar_demux_081:sink_endofpacket
	wire          id_router_081_src_valid;                                                                          // id_router_081:src_valid -> rsp_xbar_demux_081:sink_valid
	wire          id_router_081_src_startofpacket;                                                                  // id_router_081:src_startofpacket -> rsp_xbar_demux_081:sink_startofpacket
	wire  [102:0] id_router_081_src_data;                                                                           // id_router_081:src_data -> rsp_xbar_demux_081:sink_data
	wire   [98:0] id_router_081_src_channel;                                                                        // id_router_081:src_channel -> rsp_xbar_demux_081:sink_channel
	wire          id_router_081_src_ready;                                                                          // rsp_xbar_demux_081:sink_ready -> id_router_081:src_ready
	wire          cmd_xbar_demux_001_src82_ready;                                                                   // CH4_TIMER_RST_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src82_ready
	wire          id_router_082_src_endofpacket;                                                                    // id_router_082:src_endofpacket -> rsp_xbar_demux_082:sink_endofpacket
	wire          id_router_082_src_valid;                                                                          // id_router_082:src_valid -> rsp_xbar_demux_082:sink_valid
	wire          id_router_082_src_startofpacket;                                                                  // id_router_082:src_startofpacket -> rsp_xbar_demux_082:sink_startofpacket
	wire  [102:0] id_router_082_src_data;                                                                           // id_router_082:src_data -> rsp_xbar_demux_082:sink_data
	wire   [98:0] id_router_082_src_channel;                                                                        // id_router_082:src_channel -> rsp_xbar_demux_082:sink_channel
	wire          id_router_082_src_ready;                                                                          // rsp_xbar_demux_082:sink_ready -> id_router_082:src_ready
	wire          cmd_xbar_demux_001_src83_ready;                                                                   // CH4_THRESH_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src83_ready
	wire          id_router_083_src_endofpacket;                                                                    // id_router_083:src_endofpacket -> rsp_xbar_demux_083:sink_endofpacket
	wire          id_router_083_src_valid;                                                                          // id_router_083:src_valid -> rsp_xbar_demux_083:sink_valid
	wire          id_router_083_src_startofpacket;                                                                  // id_router_083:src_startofpacket -> rsp_xbar_demux_083:sink_startofpacket
	wire  [102:0] id_router_083_src_data;                                                                           // id_router_083:src_data -> rsp_xbar_demux_083:sink_data
	wire   [98:0] id_router_083_src_channel;                                                                        // id_router_083:src_channel -> rsp_xbar_demux_083:sink_channel
	wire          id_router_083_src_ready;                                                                          // rsp_xbar_demux_083:sink_ready -> id_router_083:src_ready
	wire          cmd_xbar_demux_001_src84_ready;                                                                   // CH4_RD_PEAK_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src84_ready
	wire          id_router_084_src_endofpacket;                                                                    // id_router_084:src_endofpacket -> rsp_xbar_demux_084:sink_endofpacket
	wire          id_router_084_src_valid;                                                                          // id_router_084:src_valid -> rsp_xbar_demux_084:sink_valid
	wire          id_router_084_src_startofpacket;                                                                  // id_router_084:src_startofpacket -> rsp_xbar_demux_084:sink_startofpacket
	wire  [102:0] id_router_084_src_data;                                                                           // id_router_084:src_data -> rsp_xbar_demux_084:sink_data
	wire   [98:0] id_router_084_src_channel;                                                                        // id_router_084:src_channel -> rsp_xbar_demux_084:sink_channel
	wire          id_router_084_src_ready;                                                                          // rsp_xbar_demux_084:sink_ready -> id_router_084:src_ready
	wire          cmd_xbar_demux_001_src85_ready;                                                                   // CH4_PEAK_FOUND_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src85_ready
	wire          id_router_085_src_endofpacket;                                                                    // id_router_085:src_endofpacket -> rsp_xbar_demux_085:sink_endofpacket
	wire          id_router_085_src_valid;                                                                          // id_router_085:src_valid -> rsp_xbar_demux_085:sink_valid
	wire          id_router_085_src_startofpacket;                                                                  // id_router_085:src_startofpacket -> rsp_xbar_demux_085:sink_startofpacket
	wire  [102:0] id_router_085_src_data;                                                                           // id_router_085:src_data -> rsp_xbar_demux_085:sink_data
	wire   [98:0] id_router_085_src_channel;                                                                        // id_router_085:src_channel -> rsp_xbar_demux_085:sink_channel
	wire          id_router_085_src_ready;                                                                          // rsp_xbar_demux_085:sink_ready -> id_router_085:src_ready
	wire          cmd_xbar_demux_001_src86_ready;                                                                   // CH4_TIME_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src86_ready
	wire          id_router_086_src_endofpacket;                                                                    // id_router_086:src_endofpacket -> rsp_xbar_demux_086:sink_endofpacket
	wire          id_router_086_src_valid;                                                                          // id_router_086:src_valid -> rsp_xbar_demux_086:sink_valid
	wire          id_router_086_src_startofpacket;                                                                  // id_router_086:src_startofpacket -> rsp_xbar_demux_086:sink_startofpacket
	wire  [102:0] id_router_086_src_data;                                                                           // id_router_086:src_data -> rsp_xbar_demux_086:sink_data
	wire   [98:0] id_router_086_src_channel;                                                                        // id_router_086:src_channel -> rsp_xbar_demux_086:sink_channel
	wire          id_router_086_src_ready;                                                                          // rsp_xbar_demux_086:sink_ready -> id_router_086:src_ready
	wire          cmd_xbar_demux_001_src87_ready;                                                                   // CH4_YN1_U_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src87_ready
	wire          id_router_087_src_endofpacket;                                                                    // id_router_087:src_endofpacket -> rsp_xbar_demux_087:sink_endofpacket
	wire          id_router_087_src_valid;                                                                          // id_router_087:src_valid -> rsp_xbar_demux_087:sink_valid
	wire          id_router_087_src_startofpacket;                                                                  // id_router_087:src_startofpacket -> rsp_xbar_demux_087:sink_startofpacket
	wire  [102:0] id_router_087_src_data;                                                                           // id_router_087:src_data -> rsp_xbar_demux_087:sink_data
	wire   [98:0] id_router_087_src_channel;                                                                        // id_router_087:src_channel -> rsp_xbar_demux_087:sink_channel
	wire          id_router_087_src_ready;                                                                          // rsp_xbar_demux_087:sink_ready -> id_router_087:src_ready
	wire          cmd_xbar_demux_001_src88_ready;                                                                   // CH4_YN1_MU_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src88_ready
	wire          id_router_088_src_endofpacket;                                                                    // id_router_088:src_endofpacket -> rsp_xbar_demux_088:sink_endofpacket
	wire          id_router_088_src_valid;                                                                          // id_router_088:src_valid -> rsp_xbar_demux_088:sink_valid
	wire          id_router_088_src_startofpacket;                                                                  // id_router_088:src_startofpacket -> rsp_xbar_demux_088:sink_startofpacket
	wire  [102:0] id_router_088_src_data;                                                                           // id_router_088:src_data -> rsp_xbar_demux_088:sink_data
	wire   [98:0] id_router_088_src_channel;                                                                        // id_router_088:src_channel -> rsp_xbar_demux_088:sink_channel
	wire          id_router_088_src_ready;                                                                          // rsp_xbar_demux_088:sink_ready -> id_router_088:src_ready
	wire          cmd_xbar_demux_001_src89_ready;                                                                   // CH4_YN1_ML_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src89_ready
	wire          id_router_089_src_endofpacket;                                                                    // id_router_089:src_endofpacket -> rsp_xbar_demux_089:sink_endofpacket
	wire          id_router_089_src_valid;                                                                          // id_router_089:src_valid -> rsp_xbar_demux_089:sink_valid
	wire          id_router_089_src_startofpacket;                                                                  // id_router_089:src_startofpacket -> rsp_xbar_demux_089:sink_startofpacket
	wire  [102:0] id_router_089_src_data;                                                                           // id_router_089:src_data -> rsp_xbar_demux_089:sink_data
	wire   [98:0] id_router_089_src_channel;                                                                        // id_router_089:src_channel -> rsp_xbar_demux_089:sink_channel
	wire          id_router_089_src_ready;                                                                          // rsp_xbar_demux_089:sink_ready -> id_router_089:src_ready
	wire          cmd_xbar_demux_001_src90_ready;                                                                   // CH4_YN1_L_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src90_ready
	wire          id_router_090_src_endofpacket;                                                                    // id_router_090:src_endofpacket -> rsp_xbar_demux_090:sink_endofpacket
	wire          id_router_090_src_valid;                                                                          // id_router_090:src_valid -> rsp_xbar_demux_090:sink_valid
	wire          id_router_090_src_startofpacket;                                                                  // id_router_090:src_startofpacket -> rsp_xbar_demux_090:sink_startofpacket
	wire  [102:0] id_router_090_src_data;                                                                           // id_router_090:src_data -> rsp_xbar_demux_090:sink_data
	wire   [98:0] id_router_090_src_channel;                                                                        // id_router_090:src_channel -> rsp_xbar_demux_090:sink_channel
	wire          id_router_090_src_ready;                                                                          // rsp_xbar_demux_090:sink_ready -> id_router_090:src_ready
	wire          cmd_xbar_demux_001_src91_ready;                                                                   // CH4_YN2_U_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src91_ready
	wire          id_router_091_src_endofpacket;                                                                    // id_router_091:src_endofpacket -> rsp_xbar_demux_091:sink_endofpacket
	wire          id_router_091_src_valid;                                                                          // id_router_091:src_valid -> rsp_xbar_demux_091:sink_valid
	wire          id_router_091_src_startofpacket;                                                                  // id_router_091:src_startofpacket -> rsp_xbar_demux_091:sink_startofpacket
	wire  [102:0] id_router_091_src_data;                                                                           // id_router_091:src_data -> rsp_xbar_demux_091:sink_data
	wire   [98:0] id_router_091_src_channel;                                                                        // id_router_091:src_channel -> rsp_xbar_demux_091:sink_channel
	wire          id_router_091_src_ready;                                                                          // rsp_xbar_demux_091:sink_ready -> id_router_091:src_ready
	wire          cmd_xbar_demux_001_src92_ready;                                                                   // CH4_YN2_MU_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src92_ready
	wire          id_router_092_src_endofpacket;                                                                    // id_router_092:src_endofpacket -> rsp_xbar_demux_092:sink_endofpacket
	wire          id_router_092_src_valid;                                                                          // id_router_092:src_valid -> rsp_xbar_demux_092:sink_valid
	wire          id_router_092_src_startofpacket;                                                                  // id_router_092:src_startofpacket -> rsp_xbar_demux_092:sink_startofpacket
	wire  [102:0] id_router_092_src_data;                                                                           // id_router_092:src_data -> rsp_xbar_demux_092:sink_data
	wire   [98:0] id_router_092_src_channel;                                                                        // id_router_092:src_channel -> rsp_xbar_demux_092:sink_channel
	wire          id_router_092_src_ready;                                                                          // rsp_xbar_demux_092:sink_ready -> id_router_092:src_ready
	wire          cmd_xbar_demux_001_src93_ready;                                                                   // CH4_YN2_ML_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src93_ready
	wire          id_router_093_src_endofpacket;                                                                    // id_router_093:src_endofpacket -> rsp_xbar_demux_093:sink_endofpacket
	wire          id_router_093_src_valid;                                                                          // id_router_093:src_valid -> rsp_xbar_demux_093:sink_valid
	wire          id_router_093_src_startofpacket;                                                                  // id_router_093:src_startofpacket -> rsp_xbar_demux_093:sink_startofpacket
	wire  [102:0] id_router_093_src_data;                                                                           // id_router_093:src_data -> rsp_xbar_demux_093:sink_data
	wire   [98:0] id_router_093_src_channel;                                                                        // id_router_093:src_channel -> rsp_xbar_demux_093:sink_channel
	wire          id_router_093_src_ready;                                                                          // rsp_xbar_demux_093:sink_ready -> id_router_093:src_ready
	wire          cmd_xbar_demux_001_src94_ready;                                                                   // CH4_YN2_L_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src94_ready
	wire          id_router_094_src_endofpacket;                                                                    // id_router_094:src_endofpacket -> rsp_xbar_demux_094:sink_endofpacket
	wire          id_router_094_src_valid;                                                                          // id_router_094:src_valid -> rsp_xbar_demux_094:sink_valid
	wire          id_router_094_src_startofpacket;                                                                  // id_router_094:src_startofpacket -> rsp_xbar_demux_094:sink_startofpacket
	wire  [102:0] id_router_094_src_data;                                                                           // id_router_094:src_data -> rsp_xbar_demux_094:sink_data
	wire   [98:0] id_router_094_src_channel;                                                                        // id_router_094:src_channel -> rsp_xbar_demux_094:sink_channel
	wire          id_router_094_src_ready;                                                                          // rsp_xbar_demux_094:sink_ready -> id_router_094:src_ready
	wire          cmd_xbar_demux_001_src95_ready;                                                                   // CH4_YN3_U_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src95_ready
	wire          id_router_095_src_endofpacket;                                                                    // id_router_095:src_endofpacket -> rsp_xbar_demux_095:sink_endofpacket
	wire          id_router_095_src_valid;                                                                          // id_router_095:src_valid -> rsp_xbar_demux_095:sink_valid
	wire          id_router_095_src_startofpacket;                                                                  // id_router_095:src_startofpacket -> rsp_xbar_demux_095:sink_startofpacket
	wire  [102:0] id_router_095_src_data;                                                                           // id_router_095:src_data -> rsp_xbar_demux_095:sink_data
	wire   [98:0] id_router_095_src_channel;                                                                        // id_router_095:src_channel -> rsp_xbar_demux_095:sink_channel
	wire          id_router_095_src_ready;                                                                          // rsp_xbar_demux_095:sink_ready -> id_router_095:src_ready
	wire          cmd_xbar_demux_001_src96_ready;                                                                   // CH4_YN3_MU_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src96_ready
	wire          id_router_096_src_endofpacket;                                                                    // id_router_096:src_endofpacket -> rsp_xbar_demux_096:sink_endofpacket
	wire          id_router_096_src_valid;                                                                          // id_router_096:src_valid -> rsp_xbar_demux_096:sink_valid
	wire          id_router_096_src_startofpacket;                                                                  // id_router_096:src_startofpacket -> rsp_xbar_demux_096:sink_startofpacket
	wire  [102:0] id_router_096_src_data;                                                                           // id_router_096:src_data -> rsp_xbar_demux_096:sink_data
	wire   [98:0] id_router_096_src_channel;                                                                        // id_router_096:src_channel -> rsp_xbar_demux_096:sink_channel
	wire          id_router_096_src_ready;                                                                          // rsp_xbar_demux_096:sink_ready -> id_router_096:src_ready
	wire          cmd_xbar_demux_001_src97_ready;                                                                   // CH4_YN3_ML_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src97_ready
	wire          id_router_097_src_endofpacket;                                                                    // id_router_097:src_endofpacket -> rsp_xbar_demux_097:sink_endofpacket
	wire          id_router_097_src_valid;                                                                          // id_router_097:src_valid -> rsp_xbar_demux_097:sink_valid
	wire          id_router_097_src_startofpacket;                                                                  // id_router_097:src_startofpacket -> rsp_xbar_demux_097:sink_startofpacket
	wire  [102:0] id_router_097_src_data;                                                                           // id_router_097:src_data -> rsp_xbar_demux_097:sink_data
	wire   [98:0] id_router_097_src_channel;                                                                        // id_router_097:src_channel -> rsp_xbar_demux_097:sink_channel
	wire          id_router_097_src_ready;                                                                          // rsp_xbar_demux_097:sink_ready -> id_router_097:src_ready
	wire          cmd_xbar_demux_001_src98_ready;                                                                   // CH4_YN3_L_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src98_ready
	wire          id_router_098_src_endofpacket;                                                                    // id_router_098:src_endofpacket -> rsp_xbar_demux_098:sink_endofpacket
	wire          id_router_098_src_valid;                                                                          // id_router_098:src_valid -> rsp_xbar_demux_098:sink_valid
	wire          id_router_098_src_startofpacket;                                                                  // id_router_098:src_startofpacket -> rsp_xbar_demux_098:sink_startofpacket
	wire  [102:0] id_router_098_src_data;                                                                           // id_router_098:src_data -> rsp_xbar_demux_098:sink_data
	wire   [98:0] id_router_098_src_channel;                                                                        // id_router_098:src_channel -> rsp_xbar_demux_098:sink_channel
	wire          id_router_098_src_ready;                                                                          // rsp_xbar_demux_098:sink_ready -> id_router_098:src_ready
	wire          irq_mapper_receiver0_irq;                                                                         // JTAG_UART:av_irq -> irq_mapper:receiver0_irq
	wire   [31:0] nios_cpu_d_irq_irq;                                                                               // irq_mapper:sender_irq -> NIOS_CPU:d_irq

	NIOS_SYSTEMV3_NIOS_CPU nios_cpu (
		.clk                                   (clk_clk),                                                               //                       clk.clk
		.reset_n                               (~rst_controller_reset_out_reset),                                       //                   reset_n.reset_n
		.d_address                             (nios_cpu_data_master_address),                                          //               data_master.address
		.d_byteenable                          (nios_cpu_data_master_byteenable),                                       //                          .byteenable
		.d_read                                (nios_cpu_data_master_read),                                             //                          .read
		.d_readdata                            (nios_cpu_data_master_readdata),                                         //                          .readdata
		.d_waitrequest                         (nios_cpu_data_master_waitrequest),                                      //                          .waitrequest
		.d_write                               (nios_cpu_data_master_write),                                            //                          .write
		.d_writedata                           (nios_cpu_data_master_writedata),                                        //                          .writedata
		.jtag_debug_module_debugaccess_to_roms (nios_cpu_data_master_debugaccess),                                      //                          .debugaccess
		.i_address                             (nios_cpu_instruction_master_address),                                   //        instruction_master.address
		.i_read                                (nios_cpu_instruction_master_read),                                      //                          .read
		.i_readdata                            (nios_cpu_instruction_master_readdata),                                  //                          .readdata
		.i_waitrequest                         (nios_cpu_instruction_master_waitrequest),                               //                          .waitrequest
		.d_irq                                 (nios_cpu_d_irq_irq),                                                    //                     d_irq.irq
		.jtag_debug_module_resetrequest        (nios_cpu_jtag_debug_module_reset_reset),                                //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (nios_cpu_jtag_debug_module_translator_avalon_anti_slave_0_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (nios_cpu_jtag_debug_module_translator_avalon_anti_slave_0_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (nios_cpu_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (nios_cpu_jtag_debug_module_translator_avalon_anti_slave_0_read),        //                          .read
		.jtag_debug_module_readdata            (nios_cpu_jtag_debug_module_translator_avalon_anti_slave_0_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (nios_cpu_jtag_debug_module_translator_avalon_anti_slave_0_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (nios_cpu_jtag_debug_module_translator_avalon_anti_slave_0_write),       //                          .write
		.jtag_debug_module_writedata           (nios_cpu_jtag_debug_module_translator_avalon_anti_slave_0_writedata),   //                          .writedata
		.no_ci_readra                          ()                                                                       // custom_instruction_master.readra
	);

	NIOS_SYSTEMV3_RAM ram (
		.clk        (clk_clk),                                          //   clk1.clk
		.address    (ram_s1_translator_avalon_anti_slave_0_address),    //     s1.address
		.clken      (ram_s1_translator_avalon_anti_slave_0_clken),      //       .clken
		.chipselect (ram_s1_translator_avalon_anti_slave_0_chipselect), //       .chipselect
		.write      (ram_s1_translator_avalon_anti_slave_0_write),      //       .write
		.readdata   (ram_s1_translator_avalon_anti_slave_0_readdata),   //       .readdata
		.writedata  (ram_s1_translator_avalon_anti_slave_0_writedata),  //       .writedata
		.byteenable (ram_s1_translator_avalon_anti_slave_0_byteenable), //       .byteenable
		.reset      (rst_controller_001_reset_out_reset),               // reset1.reset
		.reset_req  (rst_controller_001_reset_out_reset_req)            //       .reset_req
	);

	NIOS_SYSTEMV3_JTAG_UART jtag_uart (
		.clk            (clk_clk),                                                                //               clk.clk
		.rst_n          (~rst_controller_001_reset_out_reset),                                    //             reset.reset_n
		.av_chipselect  (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_address),     //                  .address
		.av_read_n      (~jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_read),       //                  .read_n
		.av_readdata    (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata),    //                  .readdata
		.av_write_n     (~jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_write),      //                  .write_n
		.av_writedata   (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata),   //                  .writedata
		.av_waitrequest (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                                //               irq.irq
	);

	NIOS_SYSTEMV3_LCD lcd (
		.reset_n       (~rst_controller_001_reset_out_reset),                            //         reset.reset_n
		.clk           (clk_clk),                                                        //           clk.clk
		.begintransfer (lcd_control_slave_translator_avalon_anti_slave_0_begintransfer), // control_slave.begintransfer
		.read          (lcd_control_slave_translator_avalon_anti_slave_0_read),          //              .read
		.write         (lcd_control_slave_translator_avalon_anti_slave_0_write),         //              .write
		.readdata      (lcd_control_slave_translator_avalon_anti_slave_0_readdata),      //              .readdata
		.writedata     (lcd_control_slave_translator_avalon_anti_slave_0_writedata),     //              .writedata
		.address       (lcd_control_slave_translator_avalon_anti_slave_0_address),       //              .address
		.LCD_RS        (lcd_RS),                                                         //      external.export
		.LCD_RW        (lcd_RW),                                                         //              .export
		.LCD_data      (lcd_data),                                                       //              .export
		.LCD_E         (lcd_E)                                                           //              .export
	);

	NIOS_SYSTEMV3_ADC_ON adc_on (
		.clk        (clk_clk),                                             //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                 //               reset.reset_n
		.address    (adc_on_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~adc_on_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (adc_on_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (adc_on_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (adc_on_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (adc_on_export)                                        // external_connection.export
	);

	NIOS_SYSTEMV3_FIFO_ADC_DATA fifo_adc_data (
		.clk        (clk_clk),                                                    //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                        //               reset.reset_n
		.address    (fifo_adc_data_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~fifo_adc_data_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (fifo_adc_data_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (fifo_adc_data_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (fifo_adc_data_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (fifo_adc_data_export)                                        // external_connection.export
	);

	NIOS_SYSTEMV3_ADC_ON fifo_adc_data_valid (
		.clk        (clk_clk),                                                          //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                              //               reset.reset_n
		.address    (fifo_adc_data_valid_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~fifo_adc_data_valid_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (fifo_adc_data_valid_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (fifo_adc_data_valid_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (fifo_adc_data_valid_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (fifo_adc_data_valid_export)                                        // external_connection.export
	);

	NIOS_SYSTEMV3_ADC_ON fifo_rst (
		.clk        (clk_clk),                                               //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                   //               reset.reset_n
		.address    (fifo_rst_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~fifo_rst_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (fifo_rst_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (fifo_rst_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (fifo_rst_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (fifo_rst_export)                                        // external_connection.export
	);

	NIOS_SYSTEMV3_ADC_ON subtractor_on (
		.clk        (clk_clk),                                                    //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                        //               reset.reset_n
		.address    (subtractor_on_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~subtractor_on_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (subtractor_on_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (subtractor_on_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (subtractor_on_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (subtractor_on_export)                                        // external_connection.export
	);

	NIOS_SYSTEMV3_ADC_ON ch0_timer_rst (
		.clk        (clk_clk),                                                    //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                        //               reset.reset_n
		.address    (ch0_timer_rst_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~ch0_timer_rst_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (ch0_timer_rst_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (ch0_timer_rst_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (ch0_timer_rst_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (ch0_timer_rst_export)                                        // external_connection.export
	);

	NIOS_SYSTEMV3_ADC_ON detector_on (
		.clk        (clk_clk),                                                  //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                      //               reset.reset_n
		.address    (detector_on_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~detector_on_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (detector_on_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (detector_on_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (detector_on_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (detector_on_export)                                        // external_connection.export
	);

	NIOS_SYSTEMV3_MENU menu (
		.clk        (clk_clk),                                           //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),               //               reset.reset_n
		.address    (menu_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~menu_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (menu_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (menu_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (menu_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.in_port    (menu_export)                                        // external_connection.export
	);

	NIOS_SYSTEMV3_MENU menu_up (
		.clk        (clk_clk),                                              //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                  //               reset.reset_n
		.address    (menu_up_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~menu_up_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (menu_up_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (menu_up_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (menu_up_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.in_port    (menu_up_export)                                        // external_connection.export
	);

	NIOS_SYSTEMV3_MENU_DOWN menu_down (
		.clk      (clk_clk),                                              //                 clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),                  //               reset.reset_n
		.address  (menu_down_s1_translator_avalon_anti_slave_0_address),  //                  s1.address
		.readdata (menu_down_s1_translator_avalon_anti_slave_0_readdata), //                    .readdata
		.in_port  (menu_down_export)                                      // external_connection.export
	);

	NIOS_SYSTEMV3_CH0_THRESH ch0_thresh (
		.clk        (clk_clk),                                                 //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                     //               reset.reset_n
		.address    (ch0_thresh_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~ch0_thresh_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (ch0_thresh_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (ch0_thresh_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (ch0_thresh_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (ch0_thresh_export)                                        // external_connection.export
	);

	NIOS_SYSTEMV3_ADC_ON ch0_rd_peak (
		.clk        (clk_clk),                                                  //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                      //               reset.reset_n
		.address    (ch0_rd_peak_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~ch0_rd_peak_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (ch0_rd_peak_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (ch0_rd_peak_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (ch0_rd_peak_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (ch0_rd_peak_export)                                        // external_connection.export
	);

	NIOS_SYSTEMV3_MENU ch0_peak_found (
		.clk        (clk_clk),                                                     //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                         //               reset.reset_n
		.address    (ch0_peak_found_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~ch0_peak_found_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (ch0_peak_found_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (ch0_peak_found_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (ch0_peak_found_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.in_port    (ch0_peak_found_export)                                        // external_connection.export
	);

	NIOS_SYSTEMV3_CH0_YN1_U ch0_yn1_u (
		.clk        (clk_clk),                                                //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                    //               reset.reset_n
		.address    (ch0_yn1_u_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~ch0_yn1_u_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (ch0_yn1_u_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (ch0_yn1_u_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (ch0_yn1_u_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.in_port    (ch0_yn1_u_export)                                        // external_connection.export
	);

	NIOS_SYSTEMV3_CH0_YN1_MU ch0_yn1_mu (
		.clk        (clk_clk),                                                 //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                     //               reset.reset_n
		.address    (ch0_yn1_mu_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~ch0_yn1_mu_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (ch0_yn1_mu_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (ch0_yn1_mu_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (ch0_yn1_mu_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.in_port    (ch0_yn1_mu_export)                                        // external_connection.export
	);

	NIOS_SYSTEMV3_CH0_YN1_MU ch0_yn1_ml (
		.clk        (clk_clk),                                                 //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                     //               reset.reset_n
		.address    (ch0_yn1_ml_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~ch0_yn1_ml_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (ch0_yn1_ml_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (ch0_yn1_ml_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (ch0_yn1_ml_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.in_port    (ch0_yn1_ml_export)                                        // external_connection.export
	);

	NIOS_SYSTEMV3_CH0_YN1_MU ch0_yn1_l (
		.clk        (clk_clk),                                                //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                    //               reset.reset_n
		.address    (ch0_yn1_l_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~ch0_yn1_l_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (ch0_yn1_l_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (ch0_yn1_l_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (ch0_yn1_l_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.in_port    (ch0_yn1_l_export)                                        // external_connection.export
	);

	NIOS_SYSTEMV3_CH0_YN1_U ch0_time (
		.clk        (clk_clk),                                               //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                   //               reset.reset_n
		.address    (ch0_time_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~ch0_time_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (ch0_time_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (ch0_time_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (ch0_time_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.in_port    (ch0_time_export)                                        // external_connection.export
	);

	NIOS_SYSTEMV3_CH0_YN1_U ch0_yn2_u (
		.clk        (clk_clk),                                                //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                    //               reset.reset_n
		.address    (ch0_yn2_u_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~ch0_yn2_u_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (ch0_yn2_u_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (ch0_yn2_u_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (ch0_yn2_u_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.in_port    (ch0_yn2_u_export)                                        // external_connection.export
	);

	NIOS_SYSTEMV3_CH0_YN1_MU ch0_yn2_mu (
		.clk        (clk_clk),                                                 //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                     //               reset.reset_n
		.address    (ch0_yn2_mu_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~ch0_yn2_mu_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (ch0_yn2_mu_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (ch0_yn2_mu_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (ch0_yn2_mu_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.in_port    (ch0_yn2_mu_export)                                        // external_connection.export
	);

	NIOS_SYSTEMV3_CH0_YN1_MU ch0_yn2_ml (
		.clk        (clk_clk),                                                 //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                     //               reset.reset_n
		.address    (ch0_yn2_ml_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~ch0_yn2_ml_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (ch0_yn2_ml_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (ch0_yn2_ml_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (ch0_yn2_ml_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.in_port    (ch0_yn2_ml_export)                                        // external_connection.export
	);

	NIOS_SYSTEMV3_CH0_YN1_MU ch0_yn2_l (
		.clk        (clk_clk),                                                //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                    //               reset.reset_n
		.address    (ch0_yn2_l_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~ch0_yn2_l_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (ch0_yn2_l_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (ch0_yn2_l_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (ch0_yn2_l_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.in_port    (ch0_yn2_l_export)                                        // external_connection.export
	);

	NIOS_SYSTEMV3_CH0_YN1_U ch0_yn3_u (
		.clk        (clk_clk),                                                //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                    //               reset.reset_n
		.address    (ch0_yn3_u_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~ch0_yn3_u_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (ch0_yn3_u_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (ch0_yn3_u_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (ch0_yn3_u_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.in_port    (ch0_yn3_u_export)                                        // external_connection.export
	);

	NIOS_SYSTEMV3_CH0_YN1_MU ch0_yn3_mu (
		.clk        (clk_clk),                                                 //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                     //               reset.reset_n
		.address    (ch0_yn3_mu_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~ch0_yn3_mu_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (ch0_yn3_mu_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (ch0_yn3_mu_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (ch0_yn3_mu_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.in_port    (ch0_yn3_mu_export)                                        // external_connection.export
	);

	NIOS_SYSTEMV3_CH0_YN1_MU ch0_yn3_ml (
		.clk        (clk_clk),                                                 //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                     //               reset.reset_n
		.address    (ch0_yn3_ml_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~ch0_yn3_ml_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (ch0_yn3_ml_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (ch0_yn3_ml_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (ch0_yn3_ml_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.in_port    (ch0_yn3_ml_export)                                        // external_connection.export
	);

	NIOS_SYSTEMV3_CH0_YN1_MU ch0_yn3_l (
		.clk        (clk_clk),                                                //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                    //               reset.reset_n
		.address    (ch0_yn3_l_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~ch0_yn3_l_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (ch0_yn3_l_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (ch0_yn3_l_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (ch0_yn3_l_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.in_port    (ch0_yn3_l_export)                                        // external_connection.export
	);

	NIOS_SYSTEMV3_ADC_ON ch1_timer_rst (
		.clk        (clk_clk),                                                    //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                        //               reset.reset_n
		.address    (ch1_timer_rst_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~ch1_timer_rst_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (ch1_timer_rst_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (ch1_timer_rst_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (ch1_timer_rst_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (ch1_timer_rst_export)                                        // external_connection.export
	);

	NIOS_SYSTEMV3_CH0_THRESH ch1_thresh (
		.clk        (clk_clk),                                                 //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                     //               reset.reset_n
		.address    (ch1_thresh_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~ch1_thresh_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (ch1_thresh_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (ch1_thresh_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (ch1_thresh_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (ch1_thresh_export)                                        // external_connection.export
	);

	NIOS_SYSTEMV3_ADC_ON ch1_rd_peak (
		.clk        (clk_clk),                                                  //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                      //               reset.reset_n
		.address    (ch1_rd_peak_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~ch1_rd_peak_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (ch1_rd_peak_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (ch1_rd_peak_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (ch1_rd_peak_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (ch1_rd_peak_export)                                        // external_connection.export
	);

	NIOS_SYSTEMV3_MENU ch1_peak_found (
		.clk        (clk_clk),                                                     //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                         //               reset.reset_n
		.address    (ch1_peak_found_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~ch1_peak_found_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (ch1_peak_found_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (ch1_peak_found_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (ch1_peak_found_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.in_port    (ch1_peak_found_export)                                        // external_connection.export
	);

	NIOS_SYSTEMV3_CH0_YN1_U ch1_yn1_u (
		.clk        (clk_clk),                                                //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                    //               reset.reset_n
		.address    (ch1_yn1_u_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~ch1_yn1_u_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (ch1_yn1_u_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (ch1_yn1_u_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (ch1_yn1_u_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.in_port    (ch1_yn1_u_export)                                        // external_connection.export
	);

	NIOS_SYSTEMV3_CH0_YN1_MU ch1_yn1_mu (
		.clk        (clk_clk),                                                 //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                     //               reset.reset_n
		.address    (ch1_yn1_mu_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~ch1_yn1_mu_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (ch1_yn1_mu_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (ch1_yn1_mu_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (ch1_yn1_mu_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.in_port    (ch1_yn1_mu_export)                                        // external_connection.export
	);

	NIOS_SYSTEMV3_CH0_YN1_MU ch1_yn1_ml (
		.clk        (clk_clk),                                                 //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                     //               reset.reset_n
		.address    (ch1_yn1_ml_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~ch1_yn1_ml_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (ch1_yn1_ml_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (ch1_yn1_ml_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (ch1_yn1_ml_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.in_port    (ch1_yn1_ml_export)                                        // external_connection.export
	);

	NIOS_SYSTEMV3_CH0_YN1_MU ch1_yn1_l (
		.clk        (clk_clk),                                                //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                    //               reset.reset_n
		.address    (ch1_yn1_l_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~ch1_yn1_l_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (ch1_yn1_l_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (ch1_yn1_l_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (ch1_yn1_l_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.in_port    (ch1_yn1_l_export)                                        // external_connection.export
	);

	NIOS_SYSTEMV3_CH0_YN1_U ch1_yn2_u (
		.clk        (clk_clk),                                                //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                    //               reset.reset_n
		.address    (ch1_yn2_u_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~ch1_yn2_u_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (ch1_yn2_u_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (ch1_yn2_u_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (ch1_yn2_u_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.in_port    (ch1_yn2_u_export)                                        // external_connection.export
	);

	NIOS_SYSTEMV3_CH0_YN1_MU ch1_yn2_mu (
		.clk        (clk_clk),                                                 //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                     //               reset.reset_n
		.address    (ch1_yn2_mu_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~ch1_yn2_mu_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (ch1_yn2_mu_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (ch1_yn2_mu_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (ch1_yn2_mu_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.in_port    (ch1_yn2_mu_export)                                        // external_connection.export
	);

	NIOS_SYSTEMV3_CH0_YN1_MU ch1_yn2_ml (
		.clk        (clk_clk),                                                 //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                     //               reset.reset_n
		.address    (ch1_yn2_ml_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~ch1_yn2_ml_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (ch1_yn2_ml_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (ch1_yn2_ml_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (ch1_yn2_ml_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.in_port    (ch1_yn2_ml_export)                                        // external_connection.export
	);

	NIOS_SYSTEMV3_CH0_YN1_MU ch1_yn2_l (
		.clk        (clk_clk),                                                //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                    //               reset.reset_n
		.address    (ch1_yn2_l_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~ch1_yn2_l_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (ch1_yn2_l_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (ch1_yn2_l_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (ch1_yn2_l_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.in_port    (ch1_yn2_l_export)                                        // external_connection.export
	);

	NIOS_SYSTEMV3_CH0_YN1_U ch1_yn3_u (
		.clk        (clk_clk),                                                //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                    //               reset.reset_n
		.address    (ch1_yn3_u_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~ch1_yn3_u_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (ch1_yn3_u_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (ch1_yn3_u_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (ch1_yn3_u_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.in_port    (ch1_yn3_u_export)                                        // external_connection.export
	);

	NIOS_SYSTEMV3_CH0_YN1_MU ch1_yn3_mu (
		.clk        (clk_clk),                                                 //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                     //               reset.reset_n
		.address    (ch1_yn3_mu_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~ch1_yn3_mu_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (ch1_yn3_mu_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (ch1_yn3_mu_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (ch1_yn3_mu_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.in_port    (ch1_yn3_mu_export)                                        // external_connection.export
	);

	NIOS_SYSTEMV3_CH0_YN1_MU ch1_yn3_ml (
		.clk        (clk_clk),                                                 //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                     //               reset.reset_n
		.address    (ch1_yn3_ml_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~ch1_yn3_ml_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (ch1_yn3_ml_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (ch1_yn3_ml_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (ch1_yn3_ml_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.in_port    (ch1_yn3_ml_export)                                        // external_connection.export
	);

	NIOS_SYSTEMV3_CH0_YN1_MU ch1_yn3_l (
		.clk        (clk_clk),                                                //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                    //               reset.reset_n
		.address    (ch1_yn3_l_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~ch1_yn3_l_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (ch1_yn3_l_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (ch1_yn3_l_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (ch1_yn3_l_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.in_port    (ch1_yn3_l_export)                                        // external_connection.export
	);

	NIOS_SYSTEMV3_CH0_YN1_U ch1_time (
		.clk        (clk_clk),                                               //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                   //               reset.reset_n
		.address    (ch1_time_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~ch1_time_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (ch1_time_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (ch1_time_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (ch1_time_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.in_port    (ch1_time_export)                                        // external_connection.export
	);

	NIOS_SYSTEMV3_ADC_ON ch2_timer_rst (
		.clk        (clk_clk),                                                    //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                        //               reset.reset_n
		.address    (ch2_timer_rst_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~ch2_timer_rst_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (ch2_timer_rst_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (ch2_timer_rst_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (ch2_timer_rst_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (ch2_timer_rst_export)                                        // external_connection.export
	);

	NIOS_SYSTEMV3_CH0_THRESH ch2_thresh (
		.clk        (clk_clk),                                                 //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                     //               reset.reset_n
		.address    (ch2_thresh_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~ch2_thresh_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (ch2_thresh_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (ch2_thresh_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (ch2_thresh_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (ch2_thresh_export)                                        // external_connection.export
	);

	NIOS_SYSTEMV3_ADC_ON ch2_rd_peak (
		.clk        (clk_clk),                                                  //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                      //               reset.reset_n
		.address    (ch2_rd_peak_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~ch2_rd_peak_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (ch2_rd_peak_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (ch2_rd_peak_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (ch2_rd_peak_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (ch2_rd_peak_export)                                        // external_connection.export
	);

	NIOS_SYSTEMV3_MENU ch2_peak_found (
		.clk        (clk_clk),                                                     //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                         //               reset.reset_n
		.address    (ch2_peak_found_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~ch2_peak_found_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (ch2_peak_found_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (ch2_peak_found_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (ch2_peak_found_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.in_port    (ch2_peak_found_export)                                        // external_connection.export
	);

	NIOS_SYSTEMV3_CH0_YN1_U ch2_time (
		.clk        (clk_clk),                                               //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                   //               reset.reset_n
		.address    (ch2_time_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~ch2_time_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (ch2_time_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (ch2_time_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (ch2_time_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.in_port    (ch2_time_export)                                        // external_connection.export
	);

	NIOS_SYSTEMV3_CH0_YN1_U ch2_yn1_u (
		.clk        (clk_clk),                                                //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                    //               reset.reset_n
		.address    (ch2_yn1_u_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~ch2_yn1_u_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (ch2_yn1_u_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (ch2_yn1_u_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (ch2_yn1_u_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.in_port    (ch2_yn1_u_export)                                        // external_connection.export
	);

	NIOS_SYSTEMV3_CH0_YN1_MU ch2_yn1_mu (
		.clk        (clk_clk),                                                 //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                     //               reset.reset_n
		.address    (ch2_yn1_mu_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~ch2_yn1_mu_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (ch2_yn1_mu_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (ch2_yn1_mu_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (ch2_yn1_mu_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.in_port    (ch2_yn1_mu_export)                                        // external_connection.export
	);

	NIOS_SYSTEMV3_CH0_YN1_MU ch2_yn1_ml (
		.clk        (clk_clk),                                                 //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                     //               reset.reset_n
		.address    (ch2_yn1_ml_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~ch2_yn1_ml_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (ch2_yn1_ml_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (ch2_yn1_ml_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (ch2_yn1_ml_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.in_port    (ch2_yn1_ml_export)                                        // external_connection.export
	);

	NIOS_SYSTEMV3_CH0_YN1_MU ch2_yn1_l (
		.clk        (clk_clk),                                                //                 clk.clk
		.reset_n    (~nios_cpu_jtag_debug_module_reset_reset),                //               reset.reset_n
		.address    (ch2_yn1_l_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~ch2_yn1_l_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (ch2_yn1_l_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (ch2_yn1_l_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (ch2_yn1_l_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.in_port    (ch2_yn1_l_export)                                        // external_connection.export
	);

	NIOS_SYSTEMV3_CH0_YN1_U ch2_yn2_u (
		.clk        (clk_clk),                                                //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                    //               reset.reset_n
		.address    (ch2_yn2_u_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~ch2_yn2_u_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (ch2_yn2_u_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (ch2_yn2_u_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (ch2_yn2_u_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.in_port    (ch2_yn2_u_export)                                        // external_connection.export
	);

	NIOS_SYSTEMV3_CH0_YN1_MU ch2_yn2_mu (
		.clk        (clk_clk),                                                 //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                     //               reset.reset_n
		.address    (ch2_yn2_mu_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~ch2_yn2_mu_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (ch2_yn2_mu_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (ch2_yn2_mu_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (ch2_yn2_mu_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.in_port    (ch2_yn2_mu_export)                                        // external_connection.export
	);

	NIOS_SYSTEMV3_CH0_YN1_MU ch2_yn2_ml (
		.clk        (clk_clk),                                                 //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                     //               reset.reset_n
		.address    (ch2_yn2_ml_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~ch2_yn2_ml_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (ch2_yn2_ml_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (ch2_yn2_ml_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (ch2_yn2_ml_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.in_port    (ch2_yn2_ml_export)                                        // external_connection.export
	);

	NIOS_SYSTEMV3_CH0_YN1_MU ch2_yn2_l (
		.clk        (clk_clk),                                                //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                    //               reset.reset_n
		.address    (ch2_yn2_l_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~ch2_yn2_l_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (ch2_yn2_l_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (ch2_yn2_l_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (ch2_yn2_l_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.in_port    (ch2_yn2_l_export)                                        // external_connection.export
	);

	NIOS_SYSTEMV3_CH0_YN1_U ch2_yn3_u (
		.clk        (clk_clk),                                                //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                    //               reset.reset_n
		.address    (ch2_yn3_u_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~ch2_yn3_u_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (ch2_yn3_u_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (ch2_yn3_u_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (ch2_yn3_u_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.in_port    (ch2_yn3_u_export)                                        // external_connection.export
	);

	NIOS_SYSTEMV3_CH0_YN1_MU ch2_yn3_mu (
		.clk        (clk_clk),                                                 //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                     //               reset.reset_n
		.address    (ch2_yn3_mu_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~ch2_yn3_mu_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (ch2_yn3_mu_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (ch2_yn3_mu_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (ch2_yn3_mu_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.in_port    (ch2_yn3_mu_export)                                        // external_connection.export
	);

	NIOS_SYSTEMV3_CH0_YN1_MU ch2_yn3_ml (
		.clk        (clk_clk),                                                 //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                     //               reset.reset_n
		.address    (ch2_yn3_ml_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~ch2_yn3_ml_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (ch2_yn3_ml_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (ch2_yn3_ml_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (ch2_yn3_ml_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.in_port    (ch2_yn3_ml_export)                                        // external_connection.export
	);

	NIOS_SYSTEMV3_CH0_YN1_MU ch2_yn3_l (
		.clk        (clk_clk),                                                //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                    //               reset.reset_n
		.address    (ch2_yn3_l_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~ch2_yn3_l_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (ch2_yn3_l_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (ch2_yn3_l_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (ch2_yn3_l_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.in_port    (ch2_yn3_l_export)                                        // external_connection.export
	);

	NIOS_SYSTEMV3_ADC_ON ch3_timer_rst (
		.clk        (clk_clk),                                                    //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                        //               reset.reset_n
		.address    (ch3_timer_rst_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~ch3_timer_rst_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (ch3_timer_rst_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (ch3_timer_rst_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (ch3_timer_rst_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (ch3_timer_rst_export)                                        // external_connection.export
	);

	NIOS_SYSTEMV3_CH0_THRESH ch3_thresh (
		.clk        (clk_clk),                                                 //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                     //               reset.reset_n
		.address    (ch3_thresh_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~ch3_thresh_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (ch3_thresh_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (ch3_thresh_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (ch3_thresh_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (ch3_thresh_export)                                        // external_connection.export
	);

	NIOS_SYSTEMV3_ADC_ON ch3_rd_peak (
		.clk        (clk_clk),                                                  //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                      //               reset.reset_n
		.address    (ch3_rd_peak_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~ch3_rd_peak_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (ch3_rd_peak_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (ch3_rd_peak_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (ch3_rd_peak_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (ch3_rd_peak_export)                                        // external_connection.export
	);

	NIOS_SYSTEMV3_MENU ch3_peak_found (
		.clk        (clk_clk),                                                     //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                         //               reset.reset_n
		.address    (ch3_peak_found_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~ch3_peak_found_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (ch3_peak_found_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (ch3_peak_found_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (ch3_peak_found_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.in_port    (ch3_peak_found_export)                                        // external_connection.export
	);

	NIOS_SYSTEMV3_CH0_YN1_U ch3_time (
		.clk        (clk_clk),                                               //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                   //               reset.reset_n
		.address    (ch3_time_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~ch3_time_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (ch3_time_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (ch3_time_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (ch3_time_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.in_port    (ch3_time_export)                                        // external_connection.export
	);

	NIOS_SYSTEMV3_CH0_YN1_U ch3_yn1_u (
		.clk        (clk_clk),                                                //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                    //               reset.reset_n
		.address    (ch3_yn1_u_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~ch3_yn1_u_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (ch3_yn1_u_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (ch3_yn1_u_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (ch3_yn1_u_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.in_port    (ch3_yn1_u_export)                                        // external_connection.export
	);

	NIOS_SYSTEMV3_CH0_YN1_MU ch3_yn1_mu (
		.clk        (clk_clk),                                                 //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                     //               reset.reset_n
		.address    (ch3_yn1_mu_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~ch3_yn1_mu_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (ch3_yn1_mu_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (ch3_yn1_mu_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (ch3_yn1_mu_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.in_port    (ch3_yn1_mu_export)                                        // external_connection.export
	);

	NIOS_SYSTEMV3_CH0_YN1_MU ch3_yn1_ml (
		.clk        (clk_clk),                                                 //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                     //               reset.reset_n
		.address    (ch3_yn1_ml_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~ch3_yn1_ml_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (ch3_yn1_ml_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (ch3_yn1_ml_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (ch3_yn1_ml_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.in_port    (ch3_yn1_ml_export)                                        // external_connection.export
	);

	NIOS_SYSTEMV3_CH0_YN1_MU ch3_yn1_l (
		.clk        (clk_clk),                                                //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                    //               reset.reset_n
		.address    (ch3_yn1_l_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~ch3_yn1_l_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (ch3_yn1_l_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (ch3_yn1_l_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (ch3_yn1_l_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.in_port    (ch3_yn1_l_export)                                        // external_connection.export
	);

	NIOS_SYSTEMV3_CH0_YN1_U ch3_yn2_u (
		.clk        (clk_clk),                                                //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                    //               reset.reset_n
		.address    (ch3_yn2_u_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~ch3_yn2_u_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (ch3_yn2_u_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (ch3_yn2_u_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (ch3_yn2_u_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.in_port    (ch3_yn2_u_export)                                        // external_connection.export
	);

	NIOS_SYSTEMV3_CH0_YN1_MU ch3_yn2_mu (
		.clk        (clk_clk),                                                 //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                     //               reset.reset_n
		.address    (ch3_yn2_mu_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~ch3_yn2_mu_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (ch3_yn2_mu_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (ch3_yn2_mu_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (ch3_yn2_mu_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.in_port    (ch3_yn2_mu_export)                                        // external_connection.export
	);

	NIOS_SYSTEMV3_CH0_YN1_MU ch3_yn2_ml (
		.clk        (clk_clk),                                                 //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                     //               reset.reset_n
		.address    (ch3_yn2_ml_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~ch3_yn2_ml_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (ch3_yn2_ml_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (ch3_yn2_ml_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (ch3_yn2_ml_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.in_port    (ch3_yn2_ml_export)                                        // external_connection.export
	);

	NIOS_SYSTEMV3_CH0_YN1_MU ch3_yn2_l (
		.clk        (clk_clk),                                                //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                    //               reset.reset_n
		.address    (ch3_yn2_l_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~ch3_yn2_l_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (ch3_yn2_l_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (ch3_yn2_l_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (ch3_yn2_l_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.in_port    (ch3_yn2_l_export)                                        // external_connection.export
	);

	NIOS_SYSTEMV3_CH0_YN1_U ch3_yn3_u (
		.clk        (clk_clk),                                                //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                    //               reset.reset_n
		.address    (ch3_yn3_u_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~ch3_yn3_u_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (ch3_yn3_u_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (ch3_yn3_u_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (ch3_yn3_u_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.in_port    (ch3_yn3_u_export)                                        // external_connection.export
	);

	NIOS_SYSTEMV3_CH0_YN1_MU ch3_yn3_mu (
		.clk        (clk_clk),                                                 //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                     //               reset.reset_n
		.address    (ch3_yn3_mu_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~ch3_yn3_mu_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (ch3_yn3_mu_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (ch3_yn3_mu_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (ch3_yn3_mu_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.in_port    (ch3_yn3_mu_export)                                        // external_connection.export
	);

	NIOS_SYSTEMV3_CH0_YN1_MU ch3_yn3_ml (
		.clk        (clk_clk),                                                 //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                     //               reset.reset_n
		.address    (ch3_yn3_ml_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~ch3_yn3_ml_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (ch3_yn3_ml_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (ch3_yn3_ml_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (ch3_yn3_ml_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.in_port    (ch3_yn3_ml_export)                                        // external_connection.export
	);

	NIOS_SYSTEMV3_CH0_YN1_MU ch3_yn3_l (
		.clk        (clk_clk),                                                //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                    //               reset.reset_n
		.address    (ch3_yn3_l_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~ch3_yn3_l_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (ch3_yn3_l_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (ch3_yn3_l_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (ch3_yn3_l_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.in_port    (ch3_yn3_l_export)                                        // external_connection.export
	);

	NIOS_SYSTEMV3_ADC_ON ch4_timer_rst (
		.clk        (clk_clk),                                                    //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                        //               reset.reset_n
		.address    (ch4_timer_rst_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~ch4_timer_rst_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (ch4_timer_rst_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (ch4_timer_rst_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (ch4_timer_rst_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (ch4_timer_rst_export)                                        // external_connection.export
	);

	NIOS_SYSTEMV3_CH0_THRESH ch4_thresh (
		.clk        (clk_clk),                                                 //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                     //               reset.reset_n
		.address    (ch4_thresh_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~ch4_thresh_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (ch4_thresh_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (ch4_thresh_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (ch4_thresh_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (ch4_thresh_export)                                        // external_connection.export
	);

	NIOS_SYSTEMV3_ADC_ON ch4_rd_peak (
		.clk        (clk_clk),                                                  //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                      //               reset.reset_n
		.address    (ch4_rd_peak_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~ch4_rd_peak_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (ch4_rd_peak_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (ch4_rd_peak_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (ch4_rd_peak_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (ch4_rd_peak_export)                                        // external_connection.export
	);

	NIOS_SYSTEMV3_MENU ch4_peak_found (
		.clk        (clk_clk),                                                     //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                         //               reset.reset_n
		.address    (ch4_peak_found_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~ch4_peak_found_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (ch4_peak_found_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (ch4_peak_found_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (ch4_peak_found_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.in_port    (ch4_peak_found_export)                                        // external_connection.export
	);

	NIOS_SYSTEMV3_CH0_YN1_U ch4_time (
		.clk        (clk_clk),                                               //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                   //               reset.reset_n
		.address    (ch4_time_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~ch4_time_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (ch4_time_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (ch4_time_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (ch4_time_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.in_port    (ch4_time_export)                                        // external_connection.export
	);

	NIOS_SYSTEMV3_CH0_YN1_U ch4_yn1_u (
		.clk        (clk_clk),                                                //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                    //               reset.reset_n
		.address    (ch4_yn1_u_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~ch4_yn1_u_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (ch4_yn1_u_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (ch4_yn1_u_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (ch4_yn1_u_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.in_port    (ch4_yn1_u_export)                                        // external_connection.export
	);

	NIOS_SYSTEMV3_CH0_YN1_MU ch4_yn1_mu (
		.clk        (clk_clk),                                                 //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                     //               reset.reset_n
		.address    (ch4_yn1_mu_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~ch4_yn1_mu_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (ch4_yn1_mu_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (ch4_yn1_mu_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (ch4_yn1_mu_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.in_port    (ch4_yn1_mu_export)                                        // external_connection.export
	);

	NIOS_SYSTEMV3_CH0_YN1_MU ch4_yn1_ml (
		.clk        (clk_clk),                                                 //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                     //               reset.reset_n
		.address    (ch4_yn1_ml_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~ch4_yn1_ml_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (ch4_yn1_ml_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (ch4_yn1_ml_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (ch4_yn1_ml_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.in_port    (ch4_yn1_ml_export)                                        // external_connection.export
	);

	NIOS_SYSTEMV3_CH0_YN1_MU ch4_yn1_l (
		.clk        (clk_clk),                                                //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                    //               reset.reset_n
		.address    (ch4_yn1_l_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~ch4_yn1_l_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (ch4_yn1_l_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (ch4_yn1_l_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (ch4_yn1_l_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.in_port    (ch4_yn1_l_export)                                        // external_connection.export
	);

	NIOS_SYSTEMV3_CH0_YN1_U ch4_yn2_u (
		.clk        (clk_clk),                                                //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                    //               reset.reset_n
		.address    (ch4_yn2_u_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~ch4_yn2_u_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (ch4_yn2_u_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (ch4_yn2_u_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (ch4_yn2_u_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.in_port    (ch4_yn2_u_export)                                        // external_connection.export
	);

	NIOS_SYSTEMV3_CH0_YN1_MU ch4_yn2_mu (
		.clk        (clk_clk),                                                 //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                     //               reset.reset_n
		.address    (ch4_yn2_mu_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~ch4_yn2_mu_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (ch4_yn2_mu_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (ch4_yn2_mu_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (ch4_yn2_mu_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.in_port    (ch4_yn2_mu_export)                                        // external_connection.export
	);

	NIOS_SYSTEMV3_CH0_YN1_MU ch4_yn2_ml (
		.clk        (clk_clk),                                                 //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                     //               reset.reset_n
		.address    (ch4_yn2_ml_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~ch4_yn2_ml_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (ch4_yn2_ml_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (ch4_yn2_ml_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (ch4_yn2_ml_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.in_port    (ch4_yn2_ml_export)                                        // external_connection.export
	);

	NIOS_SYSTEMV3_CH0_YN1_MU ch4_yn2_l (
		.clk        (clk_clk),                                                //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                    //               reset.reset_n
		.address    (ch4_yn2_l_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~ch4_yn2_l_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (ch4_yn2_l_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (ch4_yn2_l_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (ch4_yn2_l_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.in_port    (ch4_yn2_l_export)                                        // external_connection.export
	);

	NIOS_SYSTEMV3_CH0_YN1_U ch4_yn3_u (
		.clk        (clk_clk),                                                //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                    //               reset.reset_n
		.address    (ch4_yn3_u_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~ch4_yn3_u_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (ch4_yn3_u_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (ch4_yn3_u_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (ch4_yn3_u_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.in_port    (ch4_yn3_u_export)                                        // external_connection.export
	);

	NIOS_SYSTEMV3_CH0_YN1_MU ch4_yn3_mu (
		.clk        (clk_clk),                                                 //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                     //               reset.reset_n
		.address    (ch4_yn3_mu_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~ch4_yn3_mu_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (ch4_yn3_mu_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (ch4_yn3_mu_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (ch4_yn3_mu_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.in_port    (ch4_yn3_mu_export)                                        // external_connection.export
	);

	NIOS_SYSTEMV3_CH0_YN1_MU ch4_yn3_ml (
		.clk        (clk_clk),                                                 //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                     //               reset.reset_n
		.address    (ch4_yn3_ml_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~ch4_yn3_ml_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (ch4_yn3_ml_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (ch4_yn3_ml_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (ch4_yn3_ml_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.in_port    (ch4_yn3_ml_export)                                        // external_connection.export
	);

	NIOS_SYSTEMV3_CH0_YN1_MU ch4_yn3_l (
		.clk        (clk_clk),                                                //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                    //               reset.reset_n
		.address    (ch4_yn3_l_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~ch4_yn3_l_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (ch4_yn3_l_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (ch4_yn3_l_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (ch4_yn3_l_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.in_port    (ch4_yn3_l_export)                                        // external_connection.export
	);

	NIOS_SYSTEMV3_SSRAM #(
		.TCM_ADDRESS_W                  (21),
		.TCM_DATA_W                     (32),
		.TCM_BYTEENABLE_W               (4),
		.TCM_READ_WAIT                  (0),
		.TCM_WRITE_WAIT                 (0),
		.TCM_SETUP_WAIT                 (0),
		.TCM_DATA_HOLD                  (0),
		.TCM_TURNAROUND_TIME            (2),
		.TCM_TIMING_UNITS               (1),
		.TCM_READLATENCY                (4),
		.TCM_SYMBOLS_PER_WORD           (4),
		.USE_READDATA                   (1),
		.USE_WRITEDATA                  (1),
		.USE_READ                       (0),
		.USE_WRITE                      (1),
		.USE_BYTEENABLE                 (1),
		.USE_CHIPSELECT                 (1),
		.USE_LOCK                       (0),
		.USE_ADDRESS                    (1),
		.USE_WAITREQUEST                (0),
		.USE_WRITEBYTEENABLE            (0),
		.USE_OUTPUTENABLE               (1),
		.USE_RESETREQUEST               (0),
		.USE_IRQ                        (0),
		.USE_RESET_OUTPUT               (1),
		.ACTIVE_LOW_READ                (0),
		.ACTIVE_LOW_LOCK                (0),
		.ACTIVE_LOW_WRITE               (1),
		.ACTIVE_LOW_CHIPSELECT          (1),
		.ACTIVE_LOW_BYTEENABLE          (1),
		.ACTIVE_LOW_OUTPUTENABLE        (1),
		.ACTIVE_LOW_WRITEBYTEENABLE     (0),
		.ACTIVE_LOW_WAITREQUEST         (0),
		.ACTIVE_LOW_BEGINTRANSFER       (1),
		.CHIPSELECT_THROUGH_READLATENCY (1)
	) ssram (
		.clk_clk                 (clk_clk),                                                //   clk.clk
		.reset_reset             (rst_controller_001_reset_out_reset),                     // reset.reset
		.uas_address             (ssram_uas_translator_avalon_anti_slave_0_address),       //   uas.address
		.uas_burstcount          (ssram_uas_translator_avalon_anti_slave_0_burstcount),    //      .burstcount
		.uas_read                (ssram_uas_translator_avalon_anti_slave_0_read),          //      .read
		.uas_write               (ssram_uas_translator_avalon_anti_slave_0_write),         //      .write
		.uas_waitrequest         (ssram_uas_translator_avalon_anti_slave_0_waitrequest),   //      .waitrequest
		.uas_readdatavalid       (ssram_uas_translator_avalon_anti_slave_0_readdatavalid), //      .readdatavalid
		.uas_byteenable          (ssram_uas_translator_avalon_anti_slave_0_byteenable),    //      .byteenable
		.uas_readdata            (ssram_uas_translator_avalon_anti_slave_0_readdata),      //      .readdata
		.uas_writedata           (ssram_uas_translator_avalon_anti_slave_0_writedata),     //      .writedata
		.uas_lock                (ssram_uas_translator_avalon_anti_slave_0_lock),          //      .lock
		.uas_debugaccess         (ssram_uas_translator_avalon_anti_slave_0_debugaccess),   //      .debugaccess
		.tcm_write_n_out         (ssram_tcm_write_n_out),                                  //   tcm.write_n_out
		.tcm_begintransfer_n_out (ssram_tcm_begintransfer_n_out),                          //      .begintransfer_n_out
		.tcm_chipselect_n_out    (ssram_tcm_chipselect_n_out),                             //      .chipselect_n_out
		.tcm_outputenable_n_out  (ssram_tcm_outputenable_n_out),                           //      .outputenable_n_out
		.tcm_reset_n_out         (ssram_tcm_reset_n_out),                                  //      .reset_n_out
		.tcm_request             (ssram_tcm_request),                                      //      .request
		.tcm_grant               (ssram_tcm_grant),                                        //      .grant
		.tcm_address_out         (ssram_tcm_address_out),                                  //      .address_out
		.tcm_byteenable_n_out    (ssram_tcm_byteenable_n_out),                             //      .byteenable_n_out
		.tcm_data_out            (ssram_tcm_data_out),                                     //      .data_out
		.tcm_data_outen          (ssram_tcm_data_outen),                                   //      .data_outen
		.tcm_data_in             (ssram_tcm_data_in)                                       //      .data_in
	);

	NIOS_SYSTEMV3_tristate_bridge_ssram_pinSharer tristate_bridge_ssram_pinsharer (
		.clk_clk                          (clk_clk),                                                              //   clk.clk
		.reset_reset                      (rst_controller_001_reset_out_reset),                                   // reset.reset
		.request                          (tristate_bridge_ssram_pinsharer_tcm_request),                          //   tcm.request
		.grant                            (tristate_bridge_ssram_pinsharer_tcm_grant),                            //      .grant
		.chipenable1_n_to_the_ssram       (tristate_bridge_ssram_pinsharer_tcm_chipenable1_n_to_the_ssram_out),   //      .chipenable1_n_to_the_ssram_out
		.bw_n_to_the_ssram                (tristate_bridge_ssram_pinsharer_tcm_bw_n_to_the_ssram_out),            //      .bw_n_to_the_ssram_out
		.outputenable_n_to_the_ssram      (tristate_bridge_ssram_pinsharer_tcm_outputenable_n_to_the_ssram_out),  //      .outputenable_n_to_the_ssram_out
		.bwe_n_to_the_ssram               (tristate_bridge_ssram_pinsharer_tcm_bwe_n_to_the_ssram_out),           //      .bwe_n_to_the_ssram_out
		.data_to_and_from_the_ssram       (tristate_bridge_ssram_pinsharer_tcm_data_to_and_from_the_ssram_out),   //      .data_to_and_from_the_ssram_out
		.data_to_and_from_the_ssram_in    (tristate_bridge_ssram_pinsharer_tcm_data_to_and_from_the_ssram_in),    //      .data_to_and_from_the_ssram_in
		.data_to_and_from_the_ssram_outen (tristate_bridge_ssram_pinsharer_tcm_data_to_and_from_the_ssram_outen), //      .data_to_and_from_the_ssram_outen
		.address_to_the_ssram             (tristate_bridge_ssram_pinsharer_tcm_address_to_the_ssram_out),         //      .address_to_the_ssram_out
		.reset_n_to_the_ssram             (tristate_bridge_ssram_pinsharer_tcm_reset_n_to_the_ssram_out),         //      .reset_n_to_the_ssram_out
		.adsc_n_to_the_ssram              (tristate_bridge_ssram_pinsharer_tcm_adsc_n_to_the_ssram_out),          //      .adsc_n_to_the_ssram_out
		.tcs0_request                     (ssram_tcm_request),                                                    //  tcs0.request
		.tcs0_grant                       (ssram_tcm_grant),                                                      //      .grant
		.tcs0_chipselect_n_out            (ssram_tcm_chipselect_n_out),                                           //      .chipselect_n_out
		.tcs0_byteenable_n_out            (ssram_tcm_byteenable_n_out),                                           //      .byteenable_n_out
		.tcs0_outputenable_n_out          (ssram_tcm_outputenable_n_out),                                         //      .outputenable_n_out
		.tcs0_write_n_out                 (ssram_tcm_write_n_out),                                                //      .write_n_out
		.tcs0_data_out                    (ssram_tcm_data_out),                                                   //      .data_out
		.tcs0_data_in                     (ssram_tcm_data_in),                                                    //      .data_in
		.tcs0_data_outen                  (ssram_tcm_data_outen),                                                 //      .data_outen
		.tcs0_address_out                 (ssram_tcm_address_out),                                                //      .address_out
		.tcs0_reset_n_out                 (ssram_tcm_reset_n_out),                                                //      .reset_n_out
		.tcs0_begintransfer_n_out         (ssram_tcm_begintransfer_n_out)                                         //      .begintransfer_n_out
	);

	NIOS_SYSTEMV3_tristate_bridge_ssram tristate_bridge_ssram (
		.clk                                  (clk_clk),                                                              //   clk.clk
		.reset                                (rst_controller_001_reset_out_reset),                                   // reset.reset
		.request                              (tristate_bridge_ssram_pinsharer_tcm_request),                          //   tcs.request
		.grant                                (tristate_bridge_ssram_pinsharer_tcm_grant),                            //      .grant
		.tcs_bwe_n_to_the_ssram               (tristate_bridge_ssram_pinsharer_tcm_bwe_n_to_the_ssram_out),           //      .bwe_n_to_the_ssram_out
		.tcs_reset_n_to_the_ssram             (tristate_bridge_ssram_pinsharer_tcm_reset_n_to_the_ssram_out),         //      .reset_n_to_the_ssram_out
		.tcs_chipenable1_n_to_the_ssram       (tristate_bridge_ssram_pinsharer_tcm_chipenable1_n_to_the_ssram_out),   //      .chipenable1_n_to_the_ssram_out
		.tcs_bw_n_to_the_ssram                (tristate_bridge_ssram_pinsharer_tcm_bw_n_to_the_ssram_out),            //      .bw_n_to_the_ssram_out
		.tcs_outputenable_n_to_the_ssram      (tristate_bridge_ssram_pinsharer_tcm_outputenable_n_to_the_ssram_out),  //      .outputenable_n_to_the_ssram_out
		.tcs_adsc_n_to_the_ssram              (tristate_bridge_ssram_pinsharer_tcm_adsc_n_to_the_ssram_out),          //      .adsc_n_to_the_ssram_out
		.tcs_address_to_the_ssram             (tristate_bridge_ssram_pinsharer_tcm_address_to_the_ssram_out),         //      .address_to_the_ssram_out
		.tcs_data_to_and_from_the_ssram       (tristate_bridge_ssram_pinsharer_tcm_data_to_and_from_the_ssram_out),   //      .data_to_and_from_the_ssram_out
		.tcs_data_to_and_from_the_ssram_outen (tristate_bridge_ssram_pinsharer_tcm_data_to_and_from_the_ssram_outen), //      .data_to_and_from_the_ssram_outen
		.tcs_data_to_and_from_the_ssram_in    (tristate_bridge_ssram_pinsharer_tcm_data_to_and_from_the_ssram_in),    //      .data_to_and_from_the_ssram_in
		.bwe_n_to_the_ssram                   (tristate_bridge_ssram_bwe_n_to_the_ssram),                             //   out.bwe_n_to_the_ssram
		.reset_n_to_the_ssram                 (tristate_bridge_ssram_reset_n_to_the_ssram),                           //      .reset_n_to_the_ssram
		.chipenable1_n_to_the_ssram           (tristate_bridge_ssram_chipenable1_n_to_the_ssram),                     //      .chipenable1_n_to_the_ssram
		.bw_n_to_the_ssram                    (tristate_bridge_ssram_bw_n_to_the_ssram),                              //      .bw_n_to_the_ssram
		.outputenable_n_to_the_ssram          (tristate_bridge_ssram_outputenable_n_to_the_ssram),                    //      .outputenable_n_to_the_ssram
		.adsc_n_to_the_ssram                  (tristate_bridge_ssram_adsc_n_to_the_ssram),                            //      .adsc_n_to_the_ssram
		.address_to_the_ssram                 (tristate_bridge_ssram_address_to_the_ssram),                           //      .address_to_the_ssram
		.data_to_and_from_the_ssram           (tristate_bridge_ssram_data_to_and_from_the_ssram)                      //      .data_to_and_from_the_ssram
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (22),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (22),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (0),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (0),
		.USE_WAITREQUEST             (1),
		.USE_READRESPONSE            (0),
		.USE_WRITERESPONSE           (0),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (1),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) nios_cpu_instruction_master_translator (
		.clk                      (clk_clk),                                                                        //                       clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                 //                     reset.reset
		.uav_address              (nios_cpu_instruction_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount           (nios_cpu_instruction_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read                 (nios_cpu_instruction_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write                (nios_cpu_instruction_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest          (nios_cpu_instruction_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid        (nios_cpu_instruction_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable           (nios_cpu_instruction_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata             (nios_cpu_instruction_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata            (nios_cpu_instruction_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock                 (nios_cpu_instruction_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess          (nios_cpu_instruction_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address               (nios_cpu_instruction_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest           (nios_cpu_instruction_master_waitrequest),                                        //                          .waitrequest
		.av_read                  (nios_cpu_instruction_master_read),                                               //                          .read
		.av_readdata              (nios_cpu_instruction_master_readdata),                                           //                          .readdata
		.av_burstcount            (1'b1),                                                                           //               (terminated)
		.av_byteenable            (4'b1111),                                                                        //               (terminated)
		.av_beginbursttransfer    (1'b0),                                                                           //               (terminated)
		.av_begintransfer         (1'b0),                                                                           //               (terminated)
		.av_chipselect            (1'b0),                                                                           //               (terminated)
		.av_readdatavalid         (),                                                                               //               (terminated)
		.av_write                 (1'b0),                                                                           //               (terminated)
		.av_writedata             (32'b00000000000000000000000000000000),                                           //               (terminated)
		.av_lock                  (1'b0),                                                                           //               (terminated)
		.av_debugaccess           (1'b0),                                                                           //               (terminated)
		.uav_clken                (),                                                                               //               (terminated)
		.av_clken                 (1'b1),                                                                           //               (terminated)
		.uav_response             (2'b00),                                                                          //               (terminated)
		.av_response              (),                                                                               //               (terminated)
		.uav_writeresponserequest (),                                                                               //               (terminated)
		.uav_writeresponsevalid   (1'b0),                                                                           //               (terminated)
		.av_writeresponserequest  (1'b0),                                                                           //               (terminated)
		.av_writeresponsevalid    ()                                                                                //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (22),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (22),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (0),
		.USE_WAITREQUEST             (1),
		.USE_READRESPONSE            (0),
		.USE_WRITERESPONSE           (0),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (1)
	) nios_cpu_data_master_translator (
		.clk                      (clk_clk),                                                                 //                       clk.clk
		.reset                    (rst_controller_reset_out_reset),                                          //                     reset.reset
		.uav_address              (nios_cpu_data_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount           (nios_cpu_data_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read                 (nios_cpu_data_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write                (nios_cpu_data_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest          (nios_cpu_data_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid        (nios_cpu_data_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable           (nios_cpu_data_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata             (nios_cpu_data_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata            (nios_cpu_data_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock                 (nios_cpu_data_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess          (nios_cpu_data_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address               (nios_cpu_data_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest           (nios_cpu_data_master_waitrequest),                                        //                          .waitrequest
		.av_byteenable            (nios_cpu_data_master_byteenable),                                         //                          .byteenable
		.av_read                  (nios_cpu_data_master_read),                                               //                          .read
		.av_readdata              (nios_cpu_data_master_readdata),                                           //                          .readdata
		.av_write                 (nios_cpu_data_master_write),                                              //                          .write
		.av_writedata             (nios_cpu_data_master_writedata),                                          //                          .writedata
		.av_debugaccess           (nios_cpu_data_master_debugaccess),                                        //                          .debugaccess
		.av_burstcount            (1'b1),                                                                    //               (terminated)
		.av_beginbursttransfer    (1'b0),                                                                    //               (terminated)
		.av_begintransfer         (1'b0),                                                                    //               (terminated)
		.av_chipselect            (1'b0),                                                                    //               (terminated)
		.av_readdatavalid         (),                                                                        //               (terminated)
		.av_lock                  (1'b0),                                                                    //               (terminated)
		.uav_clken                (),                                                                        //               (terminated)
		.av_clken                 (1'b1),                                                                    //               (terminated)
		.uav_response             (2'b00),                                                                   //               (terminated)
		.av_response              (),                                                                        //               (terminated)
		.uav_writeresponserequest (),                                                                        //               (terminated)
		.uav_writeresponsevalid   (1'b0),                                                                    //               (terminated)
		.av_writeresponserequest  (1'b0),                                                                    //               (terminated)
		.av_writeresponsevalid    ()                                                                         //               (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (9),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (22),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) nios_cpu_jtag_debug_module_translator (
		.clk                      (clk_clk),                                                                               //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                        //                    reset.reset
		.uav_address              (nios_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (nios_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (nios_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (nios_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (nios_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (nios_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (nios_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (nios_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (nios_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (nios_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (nios_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (nios_cpu_jtag_debug_module_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (nios_cpu_jtag_debug_module_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (nios_cpu_jtag_debug_module_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (nios_cpu_jtag_debug_module_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (nios_cpu_jtag_debug_module_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable            (nios_cpu_jtag_debug_module_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_waitrequest           (nios_cpu_jtag_debug_module_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_debugaccess           (nios_cpu_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess),                 //                         .debugaccess
		.av_begintransfer         (),                                                                                      //              (terminated)
		.av_beginbursttransfer    (),                                                                                      //              (terminated)
		.av_burstcount            (),                                                                                      //              (terminated)
		.av_readdatavalid         (1'b0),                                                                                  //              (terminated)
		.av_writebyteenable       (),                                                                                      //              (terminated)
		.av_lock                  (),                                                                                      //              (terminated)
		.av_chipselect            (),                                                                                      //              (terminated)
		.av_clken                 (),                                                                                      //              (terminated)
		.uav_clken                (1'b0),                                                                                  //              (terminated)
		.av_outputenable          (),                                                                                      //              (terminated)
		.uav_response             (),                                                                                      //              (terminated)
		.av_response              (2'b00),                                                                                 //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                                  //              (terminated)
		.uav_writeresponsevalid   (),                                                                                      //              (terminated)
		.av_writeresponserequest  (),                                                                                      //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                   //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (11),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (22),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ram_s1_translator (
		.clk                      (clk_clk),                                                           //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                //                    reset.reset
		.uav_address              (ram_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (ram_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (ram_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (ram_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (ram_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (ram_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (ram_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (ram_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (ram_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (ram_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (ram_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (ram_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (ram_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (ram_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (ram_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable            (ram_s1_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect            (ram_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_clken                 (ram_s1_translator_avalon_anti_slave_0_clken),                       //                         .clken
		.av_read                  (),                                                                  //              (terminated)
		.av_begintransfer         (),                                                                  //              (terminated)
		.av_beginbursttransfer    (),                                                                  //              (terminated)
		.av_burstcount            (),                                                                  //              (terminated)
		.av_readdatavalid         (1'b0),                                                              //              (terminated)
		.av_waitrequest           (1'b0),                                                              //              (terminated)
		.av_writebyteenable       (),                                                                  //              (terminated)
		.av_lock                  (),                                                                  //              (terminated)
		.uav_clken                (1'b0),                                                              //              (terminated)
		.av_debugaccess           (),                                                                  //              (terminated)
		.av_outputenable          (),                                                                  //              (terminated)
		.uav_response             (),                                                                  //              (terminated)
		.av_response              (2'b00),                                                             //              (terminated)
		.uav_writeresponserequest (1'b0),                                                              //              (terminated)
		.uav_writeresponsevalid   (),                                                                  //              (terminated)
		.av_writeresponserequest  (),                                                                  //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                               //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (21),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (3),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (22),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (1),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (1),
		.AV_BURSTCOUNT_SYMBOLS          (1),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ssram_uas_translator (
		.clk                      (clk_clk),                                                              //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                   //                    reset.reset
		.uav_address              (ssram_uas_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (ssram_uas_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (ssram_uas_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (ssram_uas_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (ssram_uas_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (ssram_uas_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (ssram_uas_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (ssram_uas_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (ssram_uas_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (ssram_uas_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (ssram_uas_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (ssram_uas_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (ssram_uas_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (ssram_uas_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (ssram_uas_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (ssram_uas_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_burstcount            (ssram_uas_translator_avalon_anti_slave_0_burstcount),                  //                         .burstcount
		.av_byteenable            (ssram_uas_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_readdatavalid         (ssram_uas_translator_avalon_anti_slave_0_readdatavalid),               //                         .readdatavalid
		.av_waitrequest           (ssram_uas_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_lock                  (ssram_uas_translator_avalon_anti_slave_0_lock),                        //                         .lock
		.av_debugaccess           (ssram_uas_translator_avalon_anti_slave_0_debugaccess),                 //                         .debugaccess
		.av_begintransfer         (),                                                                     //              (terminated)
		.av_beginbursttransfer    (),                                                                     //              (terminated)
		.av_writebyteenable       (),                                                                     //              (terminated)
		.av_chipselect            (),                                                                     //              (terminated)
		.av_clken                 (),                                                                     //              (terminated)
		.uav_clken                (1'b0),                                                                 //              (terminated)
		.av_outputenable          (),                                                                     //              (terminated)
		.uav_response             (),                                                                     //              (terminated)
		.av_response              (2'b00),                                                                //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                 //              (terminated)
		.uav_writeresponsevalid   (),                                                                     //              (terminated)
		.av_writeresponserequest  (),                                                                     //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                  //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (22),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) jtag_uart_avalon_jtag_slave_translator (
		.clk                      (clk_clk),                                                                                //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                                     //                    reset.reset
		.uav_address              (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest           (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_chipselect            (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer         (),                                                                                       //              (terminated)
		.av_beginbursttransfer    (),                                                                                       //              (terminated)
		.av_burstcount            (),                                                                                       //              (terminated)
		.av_byteenable            (),                                                                                       //              (terminated)
		.av_readdatavalid         (1'b0),                                                                                   //              (terminated)
		.av_writebyteenable       (),                                                                                       //              (terminated)
		.av_lock                  (),                                                                                       //              (terminated)
		.av_clken                 (),                                                                                       //              (terminated)
		.uav_clken                (1'b0),                                                                                   //              (terminated)
		.av_debugaccess           (),                                                                                       //              (terminated)
		.av_outputenable          (),                                                                                       //              (terminated)
		.uav_response             (),                                                                                       //              (terminated)
		.av_response              (2'b00),                                                                                  //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                                   //              (terminated)
		.uav_writeresponsevalid   (),                                                                                       //              (terminated)
		.av_writeresponserequest  (),                                                                                       //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                    //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (8),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (22),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (18),
		.AV_WRITE_WAIT_CYCLES           (18),
		.AV_SETUP_WAIT_CYCLES           (18),
		.AV_DATA_HOLD_CYCLES            (18)
	) lcd_control_slave_translator (
		.clk                      (clk_clk),                                                                      //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                           //                    reset.reset
		.uav_address              (lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (lcd_control_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (lcd_control_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (lcd_control_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (lcd_control_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (lcd_control_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_begintransfer         (lcd_control_slave_translator_avalon_anti_slave_0_begintransfer),               //                         .begintransfer
		.av_beginbursttransfer    (),                                                                             //              (terminated)
		.av_burstcount            (),                                                                             //              (terminated)
		.av_byteenable            (),                                                                             //              (terminated)
		.av_readdatavalid         (1'b0),                                                                         //              (terminated)
		.av_waitrequest           (1'b0),                                                                         //              (terminated)
		.av_writebyteenable       (),                                                                             //              (terminated)
		.av_lock                  (),                                                                             //              (terminated)
		.av_chipselect            (),                                                                             //              (terminated)
		.av_clken                 (),                                                                             //              (terminated)
		.uav_clken                (1'b0),                                                                         //              (terminated)
		.av_debugaccess           (),                                                                             //              (terminated)
		.av_outputenable          (),                                                                             //              (terminated)
		.uav_response             (),                                                                             //              (terminated)
		.av_response              (2'b00),                                                                        //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                         //              (terminated)
		.uav_writeresponsevalid   (),                                                                             //              (terminated)
		.av_writeresponserequest  (),                                                                             //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                          //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (22),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) adc_on_s1_translator (
		.clk                      (clk_clk),                                                              //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                   //                    reset.reset
		.uav_address              (adc_on_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (adc_on_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (adc_on_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (adc_on_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (adc_on_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (adc_on_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (adc_on_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (adc_on_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (adc_on_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (adc_on_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (adc_on_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (adc_on_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (adc_on_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (adc_on_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (adc_on_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (adc_on_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                     //              (terminated)
		.av_begintransfer         (),                                                                     //              (terminated)
		.av_beginbursttransfer    (),                                                                     //              (terminated)
		.av_burstcount            (),                                                                     //              (terminated)
		.av_byteenable            (),                                                                     //              (terminated)
		.av_readdatavalid         (1'b0),                                                                 //              (terminated)
		.av_waitrequest           (1'b0),                                                                 //              (terminated)
		.av_writebyteenable       (),                                                                     //              (terminated)
		.av_lock                  (),                                                                     //              (terminated)
		.av_clken                 (),                                                                     //              (terminated)
		.uav_clken                (1'b0),                                                                 //              (terminated)
		.av_debugaccess           (),                                                                     //              (terminated)
		.av_outputenable          (),                                                                     //              (terminated)
		.uav_response             (),                                                                     //              (terminated)
		.av_response              (2'b00),                                                                //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                 //              (terminated)
		.uav_writeresponsevalid   (),                                                                     //              (terminated)
		.av_writeresponserequest  (),                                                                     //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                  //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (22),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) fifo_adc_data_s1_translator (
		.clk                      (clk_clk),                                                                     //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                          //                    reset.reset
		.uav_address              (fifo_adc_data_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (fifo_adc_data_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (fifo_adc_data_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (fifo_adc_data_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (fifo_adc_data_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (fifo_adc_data_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (fifo_adc_data_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (fifo_adc_data_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (fifo_adc_data_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (fifo_adc_data_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (fifo_adc_data_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (fifo_adc_data_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (fifo_adc_data_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (fifo_adc_data_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (fifo_adc_data_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (fifo_adc_data_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                            //              (terminated)
		.av_begintransfer         (),                                                                            //              (terminated)
		.av_beginbursttransfer    (),                                                                            //              (terminated)
		.av_burstcount            (),                                                                            //              (terminated)
		.av_byteenable            (),                                                                            //              (terminated)
		.av_readdatavalid         (1'b0),                                                                        //              (terminated)
		.av_waitrequest           (1'b0),                                                                        //              (terminated)
		.av_writebyteenable       (),                                                                            //              (terminated)
		.av_lock                  (),                                                                            //              (terminated)
		.av_clken                 (),                                                                            //              (terminated)
		.uav_clken                (1'b0),                                                                        //              (terminated)
		.av_debugaccess           (),                                                                            //              (terminated)
		.av_outputenable          (),                                                                            //              (terminated)
		.uav_response             (),                                                                            //              (terminated)
		.av_response              (2'b00),                                                                       //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                        //              (terminated)
		.uav_writeresponsevalid   (),                                                                            //              (terminated)
		.av_writeresponserequest  (),                                                                            //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                         //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (22),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) fifo_adc_data_valid_s1_translator (
		.clk                      (clk_clk),                                                                           //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                                //                    reset.reset
		.uav_address              (fifo_adc_data_valid_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (fifo_adc_data_valid_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (fifo_adc_data_valid_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (fifo_adc_data_valid_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (fifo_adc_data_valid_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (fifo_adc_data_valid_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (fifo_adc_data_valid_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (fifo_adc_data_valid_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (fifo_adc_data_valid_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (fifo_adc_data_valid_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (fifo_adc_data_valid_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (fifo_adc_data_valid_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (fifo_adc_data_valid_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (fifo_adc_data_valid_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (fifo_adc_data_valid_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (fifo_adc_data_valid_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                                  //              (terminated)
		.av_begintransfer         (),                                                                                  //              (terminated)
		.av_beginbursttransfer    (),                                                                                  //              (terminated)
		.av_burstcount            (),                                                                                  //              (terminated)
		.av_byteenable            (),                                                                                  //              (terminated)
		.av_readdatavalid         (1'b0),                                                                              //              (terminated)
		.av_waitrequest           (1'b0),                                                                              //              (terminated)
		.av_writebyteenable       (),                                                                                  //              (terminated)
		.av_lock                  (),                                                                                  //              (terminated)
		.av_clken                 (),                                                                                  //              (terminated)
		.uav_clken                (1'b0),                                                                              //              (terminated)
		.av_debugaccess           (),                                                                                  //              (terminated)
		.av_outputenable          (),                                                                                  //              (terminated)
		.uav_response             (),                                                                                  //              (terminated)
		.av_response              (2'b00),                                                                             //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                              //              (terminated)
		.uav_writeresponsevalid   (),                                                                                  //              (terminated)
		.av_writeresponserequest  (),                                                                                  //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                               //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (22),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) fifo_rst_s1_translator (
		.clk                      (clk_clk),                                                                //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                     //                    reset.reset
		.uav_address              (fifo_rst_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (fifo_rst_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (fifo_rst_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (fifo_rst_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (fifo_rst_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (fifo_rst_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (fifo_rst_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (fifo_rst_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (fifo_rst_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (fifo_rst_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (fifo_rst_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (fifo_rst_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (fifo_rst_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (fifo_rst_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (fifo_rst_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (fifo_rst_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                       //              (terminated)
		.av_begintransfer         (),                                                                       //              (terminated)
		.av_beginbursttransfer    (),                                                                       //              (terminated)
		.av_burstcount            (),                                                                       //              (terminated)
		.av_byteenable            (),                                                                       //              (terminated)
		.av_readdatavalid         (1'b0),                                                                   //              (terminated)
		.av_waitrequest           (1'b0),                                                                   //              (terminated)
		.av_writebyteenable       (),                                                                       //              (terminated)
		.av_lock                  (),                                                                       //              (terminated)
		.av_clken                 (),                                                                       //              (terminated)
		.uav_clken                (1'b0),                                                                   //              (terminated)
		.av_debugaccess           (),                                                                       //              (terminated)
		.av_outputenable          (),                                                                       //              (terminated)
		.uav_response             (),                                                                       //              (terminated)
		.av_response              (2'b00),                                                                  //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                   //              (terminated)
		.uav_writeresponsevalid   (),                                                                       //              (terminated)
		.av_writeresponserequest  (),                                                                       //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                    //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (22),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) subtractor_on_s1_translator (
		.clk                      (clk_clk),                                                                     //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                          //                    reset.reset
		.uav_address              (subtractor_on_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (subtractor_on_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (subtractor_on_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (subtractor_on_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (subtractor_on_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (subtractor_on_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (subtractor_on_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (subtractor_on_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (subtractor_on_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (subtractor_on_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (subtractor_on_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (subtractor_on_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (subtractor_on_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (subtractor_on_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (subtractor_on_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (subtractor_on_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                            //              (terminated)
		.av_begintransfer         (),                                                                            //              (terminated)
		.av_beginbursttransfer    (),                                                                            //              (terminated)
		.av_burstcount            (),                                                                            //              (terminated)
		.av_byteenable            (),                                                                            //              (terminated)
		.av_readdatavalid         (1'b0),                                                                        //              (terminated)
		.av_waitrequest           (1'b0),                                                                        //              (terminated)
		.av_writebyteenable       (),                                                                            //              (terminated)
		.av_lock                  (),                                                                            //              (terminated)
		.av_clken                 (),                                                                            //              (terminated)
		.uav_clken                (1'b0),                                                                        //              (terminated)
		.av_debugaccess           (),                                                                            //              (terminated)
		.av_outputenable          (),                                                                            //              (terminated)
		.uav_response             (),                                                                            //              (terminated)
		.av_response              (2'b00),                                                                       //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                        //              (terminated)
		.uav_writeresponsevalid   (),                                                                            //              (terminated)
		.av_writeresponserequest  (),                                                                            //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                         //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (22),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ch0_timer_rst_s1_translator (
		.clk                      (clk_clk),                                                                     //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                          //                    reset.reset
		.uav_address              (ch0_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (ch0_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (ch0_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (ch0_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (ch0_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (ch0_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (ch0_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (ch0_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (ch0_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (ch0_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (ch0_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (ch0_timer_rst_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (ch0_timer_rst_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (ch0_timer_rst_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (ch0_timer_rst_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (ch0_timer_rst_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                            //              (terminated)
		.av_begintransfer         (),                                                                            //              (terminated)
		.av_beginbursttransfer    (),                                                                            //              (terminated)
		.av_burstcount            (),                                                                            //              (terminated)
		.av_byteenable            (),                                                                            //              (terminated)
		.av_readdatavalid         (1'b0),                                                                        //              (terminated)
		.av_waitrequest           (1'b0),                                                                        //              (terminated)
		.av_writebyteenable       (),                                                                            //              (terminated)
		.av_lock                  (),                                                                            //              (terminated)
		.av_clken                 (),                                                                            //              (terminated)
		.uav_clken                (1'b0),                                                                        //              (terminated)
		.av_debugaccess           (),                                                                            //              (terminated)
		.av_outputenable          (),                                                                            //              (terminated)
		.uav_response             (),                                                                            //              (terminated)
		.av_response              (2'b00),                                                                       //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                        //              (terminated)
		.uav_writeresponsevalid   (),                                                                            //              (terminated)
		.av_writeresponserequest  (),                                                                            //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                         //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (22),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) detector_on_s1_translator (
		.clk                      (clk_clk),                                                                   //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                        //                    reset.reset
		.uav_address              (detector_on_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (detector_on_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (detector_on_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (detector_on_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (detector_on_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (detector_on_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (detector_on_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (detector_on_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (detector_on_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (detector_on_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (detector_on_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (detector_on_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (detector_on_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (detector_on_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (detector_on_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (detector_on_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                          //              (terminated)
		.av_begintransfer         (),                                                                          //              (terminated)
		.av_beginbursttransfer    (),                                                                          //              (terminated)
		.av_burstcount            (),                                                                          //              (terminated)
		.av_byteenable            (),                                                                          //              (terminated)
		.av_readdatavalid         (1'b0),                                                                      //              (terminated)
		.av_waitrequest           (1'b0),                                                                      //              (terminated)
		.av_writebyteenable       (),                                                                          //              (terminated)
		.av_lock                  (),                                                                          //              (terminated)
		.av_clken                 (),                                                                          //              (terminated)
		.uav_clken                (1'b0),                                                                      //              (terminated)
		.av_debugaccess           (),                                                                          //              (terminated)
		.av_outputenable          (),                                                                          //              (terminated)
		.uav_response             (),                                                                          //              (terminated)
		.av_response              (2'b00),                                                                     //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                      //              (terminated)
		.uav_writeresponsevalid   (),                                                                          //              (terminated)
		.av_writeresponserequest  (),                                                                          //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                       //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (22),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) menu_down_s1_translator (
		.clk                      (clk_clk),                                                                 //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                      //                    reset.reset
		.uav_address              (menu_down_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (menu_down_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (menu_down_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (menu_down_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (menu_down_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (menu_down_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (menu_down_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (menu_down_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (menu_down_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (menu_down_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (menu_down_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (menu_down_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_readdata              (menu_down_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_write                 (),                                                                        //              (terminated)
		.av_read                  (),                                                                        //              (terminated)
		.av_writedata             (),                                                                        //              (terminated)
		.av_begintransfer         (),                                                                        //              (terminated)
		.av_beginbursttransfer    (),                                                                        //              (terminated)
		.av_burstcount            (),                                                                        //              (terminated)
		.av_byteenable            (),                                                                        //              (terminated)
		.av_readdatavalid         (1'b0),                                                                    //              (terminated)
		.av_waitrequest           (1'b0),                                                                    //              (terminated)
		.av_writebyteenable       (),                                                                        //              (terminated)
		.av_lock                  (),                                                                        //              (terminated)
		.av_chipselect            (),                                                                        //              (terminated)
		.av_clken                 (),                                                                        //              (terminated)
		.uav_clken                (1'b0),                                                                    //              (terminated)
		.av_debugaccess           (),                                                                        //              (terminated)
		.av_outputenable          (),                                                                        //              (terminated)
		.uav_response             (),                                                                        //              (terminated)
		.av_response              (2'b00),                                                                   //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                    //              (terminated)
		.uav_writeresponsevalid   (),                                                                        //              (terminated)
		.av_writeresponserequest  (),                                                                        //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                     //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (22),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) menu_up_s1_translator (
		.clk                      (clk_clk),                                                               //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                    //                    reset.reset
		.uav_address              (menu_up_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (menu_up_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (menu_up_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (menu_up_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (menu_up_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (menu_up_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (menu_up_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (menu_up_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (menu_up_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (menu_up_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (menu_up_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (menu_up_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (menu_up_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (menu_up_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (menu_up_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (menu_up_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                      //              (terminated)
		.av_begintransfer         (),                                                                      //              (terminated)
		.av_beginbursttransfer    (),                                                                      //              (terminated)
		.av_burstcount            (),                                                                      //              (terminated)
		.av_byteenable            (),                                                                      //              (terminated)
		.av_readdatavalid         (1'b0),                                                                  //              (terminated)
		.av_waitrequest           (1'b0),                                                                  //              (terminated)
		.av_writebyteenable       (),                                                                      //              (terminated)
		.av_lock                  (),                                                                      //              (terminated)
		.av_clken                 (),                                                                      //              (terminated)
		.uav_clken                (1'b0),                                                                  //              (terminated)
		.av_debugaccess           (),                                                                      //              (terminated)
		.av_outputenable          (),                                                                      //              (terminated)
		.uav_response             (),                                                                      //              (terminated)
		.av_response              (2'b00),                                                                 //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                  //              (terminated)
		.uav_writeresponsevalid   (),                                                                      //              (terminated)
		.av_writeresponserequest  (),                                                                      //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                   //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (22),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) menu_s1_translator (
		.clk                      (clk_clk),                                                            //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                 //                    reset.reset
		.uav_address              (menu_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (menu_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (menu_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (menu_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (menu_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (menu_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (menu_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (menu_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (menu_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (menu_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (menu_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (menu_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (menu_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (menu_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (menu_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (menu_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                   //              (terminated)
		.av_begintransfer         (),                                                                   //              (terminated)
		.av_beginbursttransfer    (),                                                                   //              (terminated)
		.av_burstcount            (),                                                                   //              (terminated)
		.av_byteenable            (),                                                                   //              (terminated)
		.av_readdatavalid         (1'b0),                                                               //              (terminated)
		.av_waitrequest           (1'b0),                                                               //              (terminated)
		.av_writebyteenable       (),                                                                   //              (terminated)
		.av_lock                  (),                                                                   //              (terminated)
		.av_clken                 (),                                                                   //              (terminated)
		.uav_clken                (1'b0),                                                               //              (terminated)
		.av_debugaccess           (),                                                                   //              (terminated)
		.av_outputenable          (),                                                                   //              (terminated)
		.uav_response             (),                                                                   //              (terminated)
		.av_response              (2'b00),                                                              //              (terminated)
		.uav_writeresponserequest (1'b0),                                                               //              (terminated)
		.uav_writeresponsevalid   (),                                                                   //              (terminated)
		.av_writeresponserequest  (),                                                                   //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (22),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ch0_thresh_s1_translator (
		.clk                      (clk_clk),                                                                  //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                       //                    reset.reset
		.uav_address              (ch0_thresh_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (ch0_thresh_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (ch0_thresh_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (ch0_thresh_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (ch0_thresh_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (ch0_thresh_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (ch0_thresh_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (ch0_thresh_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (ch0_thresh_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (ch0_thresh_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (ch0_thresh_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (ch0_thresh_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (ch0_thresh_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (ch0_thresh_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (ch0_thresh_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (ch0_thresh_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                         //              (terminated)
		.av_begintransfer         (),                                                                         //              (terminated)
		.av_beginbursttransfer    (),                                                                         //              (terminated)
		.av_burstcount            (),                                                                         //              (terminated)
		.av_byteenable            (),                                                                         //              (terminated)
		.av_readdatavalid         (1'b0),                                                                     //              (terminated)
		.av_waitrequest           (1'b0),                                                                     //              (terminated)
		.av_writebyteenable       (),                                                                         //              (terminated)
		.av_lock                  (),                                                                         //              (terminated)
		.av_clken                 (),                                                                         //              (terminated)
		.uav_clken                (1'b0),                                                                     //              (terminated)
		.av_debugaccess           (),                                                                         //              (terminated)
		.av_outputenable          (),                                                                         //              (terminated)
		.uav_response             (),                                                                         //              (terminated)
		.av_response              (2'b00),                                                                    //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                     //              (terminated)
		.uav_writeresponsevalid   (),                                                                         //              (terminated)
		.av_writeresponserequest  (),                                                                         //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                      //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (22),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ch0_rd_peak_s1_translator (
		.clk                      (clk_clk),                                                                   //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                        //                    reset.reset
		.uav_address              (ch0_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (ch0_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (ch0_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (ch0_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (ch0_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (ch0_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (ch0_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (ch0_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (ch0_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (ch0_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (ch0_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (ch0_rd_peak_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (ch0_rd_peak_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (ch0_rd_peak_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (ch0_rd_peak_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (ch0_rd_peak_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                          //              (terminated)
		.av_begintransfer         (),                                                                          //              (terminated)
		.av_beginbursttransfer    (),                                                                          //              (terminated)
		.av_burstcount            (),                                                                          //              (terminated)
		.av_byteenable            (),                                                                          //              (terminated)
		.av_readdatavalid         (1'b0),                                                                      //              (terminated)
		.av_waitrequest           (1'b0),                                                                      //              (terminated)
		.av_writebyteenable       (),                                                                          //              (terminated)
		.av_lock                  (),                                                                          //              (terminated)
		.av_clken                 (),                                                                          //              (terminated)
		.uav_clken                (1'b0),                                                                      //              (terminated)
		.av_debugaccess           (),                                                                          //              (terminated)
		.av_outputenable          (),                                                                          //              (terminated)
		.uav_response             (),                                                                          //              (terminated)
		.av_response              (2'b00),                                                                     //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                      //              (terminated)
		.uav_writeresponsevalid   (),                                                                          //              (terminated)
		.av_writeresponserequest  (),                                                                          //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                       //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (22),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ch0_peak_found_s1_translator (
		.clk                      (clk_clk),                                                                      //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                           //                    reset.reset
		.uav_address              (ch0_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (ch0_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (ch0_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (ch0_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (ch0_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (ch0_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (ch0_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (ch0_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (ch0_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (ch0_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (ch0_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (ch0_peak_found_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (ch0_peak_found_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (ch0_peak_found_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (ch0_peak_found_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (ch0_peak_found_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                             //              (terminated)
		.av_begintransfer         (),                                                                             //              (terminated)
		.av_beginbursttransfer    (),                                                                             //              (terminated)
		.av_burstcount            (),                                                                             //              (terminated)
		.av_byteenable            (),                                                                             //              (terminated)
		.av_readdatavalid         (1'b0),                                                                         //              (terminated)
		.av_waitrequest           (1'b0),                                                                         //              (terminated)
		.av_writebyteenable       (),                                                                             //              (terminated)
		.av_lock                  (),                                                                             //              (terminated)
		.av_clken                 (),                                                                             //              (terminated)
		.uav_clken                (1'b0),                                                                         //              (terminated)
		.av_debugaccess           (),                                                                             //              (terminated)
		.av_outputenable          (),                                                                             //              (terminated)
		.uav_response             (),                                                                             //              (terminated)
		.av_response              (2'b00),                                                                        //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                         //              (terminated)
		.uav_writeresponsevalid   (),                                                                             //              (terminated)
		.av_writeresponserequest  (),                                                                             //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                          //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (22),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ch0_yn1_l_s1_translator (
		.clk                      (clk_clk),                                                                 //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                      //                    reset.reset
		.uav_address              (ch0_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (ch0_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (ch0_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (ch0_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (ch0_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (ch0_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (ch0_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (ch0_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (ch0_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (ch0_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (ch0_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (ch0_yn1_l_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (ch0_yn1_l_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (ch0_yn1_l_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (ch0_yn1_l_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (ch0_yn1_l_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                        //              (terminated)
		.av_begintransfer         (),                                                                        //              (terminated)
		.av_beginbursttransfer    (),                                                                        //              (terminated)
		.av_burstcount            (),                                                                        //              (terminated)
		.av_byteenable            (),                                                                        //              (terminated)
		.av_readdatavalid         (1'b0),                                                                    //              (terminated)
		.av_waitrequest           (1'b0),                                                                    //              (terminated)
		.av_writebyteenable       (),                                                                        //              (terminated)
		.av_lock                  (),                                                                        //              (terminated)
		.av_clken                 (),                                                                        //              (terminated)
		.uav_clken                (1'b0),                                                                    //              (terminated)
		.av_debugaccess           (),                                                                        //              (terminated)
		.av_outputenable          (),                                                                        //              (terminated)
		.uav_response             (),                                                                        //              (terminated)
		.av_response              (2'b00),                                                                   //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                    //              (terminated)
		.uav_writeresponsevalid   (),                                                                        //              (terminated)
		.av_writeresponserequest  (),                                                                        //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                     //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (22),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ch0_yn1_ml_s1_translator (
		.clk                      (clk_clk),                                                                  //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                       //                    reset.reset
		.uav_address              (ch0_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (ch0_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (ch0_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (ch0_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (ch0_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (ch0_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (ch0_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (ch0_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (ch0_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (ch0_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (ch0_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (ch0_yn1_ml_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (ch0_yn1_ml_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (ch0_yn1_ml_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (ch0_yn1_ml_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (ch0_yn1_ml_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                         //              (terminated)
		.av_begintransfer         (),                                                                         //              (terminated)
		.av_beginbursttransfer    (),                                                                         //              (terminated)
		.av_burstcount            (),                                                                         //              (terminated)
		.av_byteenable            (),                                                                         //              (terminated)
		.av_readdatavalid         (1'b0),                                                                     //              (terminated)
		.av_waitrequest           (1'b0),                                                                     //              (terminated)
		.av_writebyteenable       (),                                                                         //              (terminated)
		.av_lock                  (),                                                                         //              (terminated)
		.av_clken                 (),                                                                         //              (terminated)
		.uav_clken                (1'b0),                                                                     //              (terminated)
		.av_debugaccess           (),                                                                         //              (terminated)
		.av_outputenable          (),                                                                         //              (terminated)
		.uav_response             (),                                                                         //              (terminated)
		.av_response              (2'b00),                                                                    //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                     //              (terminated)
		.uav_writeresponsevalid   (),                                                                         //              (terminated)
		.av_writeresponserequest  (),                                                                         //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                      //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (22),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ch0_yn1_mu_s1_translator (
		.clk                      (clk_clk),                                                                  //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                       //                    reset.reset
		.uav_address              (ch0_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (ch0_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (ch0_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (ch0_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (ch0_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (ch0_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (ch0_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (ch0_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (ch0_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (ch0_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (ch0_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (ch0_yn1_mu_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (ch0_yn1_mu_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (ch0_yn1_mu_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (ch0_yn1_mu_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (ch0_yn1_mu_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                         //              (terminated)
		.av_begintransfer         (),                                                                         //              (terminated)
		.av_beginbursttransfer    (),                                                                         //              (terminated)
		.av_burstcount            (),                                                                         //              (terminated)
		.av_byteenable            (),                                                                         //              (terminated)
		.av_readdatavalid         (1'b0),                                                                     //              (terminated)
		.av_waitrequest           (1'b0),                                                                     //              (terminated)
		.av_writebyteenable       (),                                                                         //              (terminated)
		.av_lock                  (),                                                                         //              (terminated)
		.av_clken                 (),                                                                         //              (terminated)
		.uav_clken                (1'b0),                                                                     //              (terminated)
		.av_debugaccess           (),                                                                         //              (terminated)
		.av_outputenable          (),                                                                         //              (terminated)
		.uav_response             (),                                                                         //              (terminated)
		.av_response              (2'b00),                                                                    //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                     //              (terminated)
		.uav_writeresponsevalid   (),                                                                         //              (terminated)
		.av_writeresponserequest  (),                                                                         //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                      //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (22),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ch0_yn1_u_s1_translator (
		.clk                      (clk_clk),                                                                 //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                      //                    reset.reset
		.uav_address              (ch0_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (ch0_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (ch0_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (ch0_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (ch0_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (ch0_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (ch0_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (ch0_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (ch0_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (ch0_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (ch0_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (ch0_yn1_u_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (ch0_yn1_u_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (ch0_yn1_u_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (ch0_yn1_u_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (ch0_yn1_u_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                        //              (terminated)
		.av_begintransfer         (),                                                                        //              (terminated)
		.av_beginbursttransfer    (),                                                                        //              (terminated)
		.av_burstcount            (),                                                                        //              (terminated)
		.av_byteenable            (),                                                                        //              (terminated)
		.av_readdatavalid         (1'b0),                                                                    //              (terminated)
		.av_waitrequest           (1'b0),                                                                    //              (terminated)
		.av_writebyteenable       (),                                                                        //              (terminated)
		.av_lock                  (),                                                                        //              (terminated)
		.av_clken                 (),                                                                        //              (terminated)
		.uav_clken                (1'b0),                                                                    //              (terminated)
		.av_debugaccess           (),                                                                        //              (terminated)
		.av_outputenable          (),                                                                        //              (terminated)
		.uav_response             (),                                                                        //              (terminated)
		.av_response              (2'b00),                                                                   //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                    //              (terminated)
		.uav_writeresponsevalid   (),                                                                        //              (terminated)
		.av_writeresponserequest  (),                                                                        //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                     //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (22),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ch0_time_s1_translator (
		.clk                      (clk_clk),                                                                //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                     //                    reset.reset
		.uav_address              (ch0_time_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (ch0_time_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (ch0_time_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (ch0_time_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (ch0_time_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (ch0_time_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (ch0_time_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (ch0_time_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (ch0_time_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (ch0_time_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (ch0_time_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (ch0_time_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (ch0_time_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (ch0_time_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (ch0_time_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (ch0_time_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                       //              (terminated)
		.av_begintransfer         (),                                                                       //              (terminated)
		.av_beginbursttransfer    (),                                                                       //              (terminated)
		.av_burstcount            (),                                                                       //              (terminated)
		.av_byteenable            (),                                                                       //              (terminated)
		.av_readdatavalid         (1'b0),                                                                   //              (terminated)
		.av_waitrequest           (1'b0),                                                                   //              (terminated)
		.av_writebyteenable       (),                                                                       //              (terminated)
		.av_lock                  (),                                                                       //              (terminated)
		.av_clken                 (),                                                                       //              (terminated)
		.uav_clken                (1'b0),                                                                   //              (terminated)
		.av_debugaccess           (),                                                                       //              (terminated)
		.av_outputenable          (),                                                                       //              (terminated)
		.uav_response             (),                                                                       //              (terminated)
		.av_response              (2'b00),                                                                  //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                   //              (terminated)
		.uav_writeresponsevalid   (),                                                                       //              (terminated)
		.av_writeresponserequest  (),                                                                       //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                    //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (22),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ch0_yn2_mu_s1_translator (
		.clk                      (clk_clk),                                                                  //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                       //                    reset.reset
		.uav_address              (ch0_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (ch0_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (ch0_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (ch0_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (ch0_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (ch0_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (ch0_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (ch0_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (ch0_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (ch0_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (ch0_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (ch0_yn2_mu_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (ch0_yn2_mu_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (ch0_yn2_mu_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (ch0_yn2_mu_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (ch0_yn2_mu_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                         //              (terminated)
		.av_begintransfer         (),                                                                         //              (terminated)
		.av_beginbursttransfer    (),                                                                         //              (terminated)
		.av_burstcount            (),                                                                         //              (terminated)
		.av_byteenable            (),                                                                         //              (terminated)
		.av_readdatavalid         (1'b0),                                                                     //              (terminated)
		.av_waitrequest           (1'b0),                                                                     //              (terminated)
		.av_writebyteenable       (),                                                                         //              (terminated)
		.av_lock                  (),                                                                         //              (terminated)
		.av_clken                 (),                                                                         //              (terminated)
		.uav_clken                (1'b0),                                                                     //              (terminated)
		.av_debugaccess           (),                                                                         //              (terminated)
		.av_outputenable          (),                                                                         //              (terminated)
		.uav_response             (),                                                                         //              (terminated)
		.av_response              (2'b00),                                                                    //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                     //              (terminated)
		.uav_writeresponsevalid   (),                                                                         //              (terminated)
		.av_writeresponserequest  (),                                                                         //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                      //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (22),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ch0_yn2_ml_s1_translator (
		.clk                      (clk_clk),                                                                  //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                       //                    reset.reset
		.uav_address              (ch0_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (ch0_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (ch0_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (ch0_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (ch0_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (ch0_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (ch0_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (ch0_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (ch0_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (ch0_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (ch0_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (ch0_yn2_ml_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (ch0_yn2_ml_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (ch0_yn2_ml_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (ch0_yn2_ml_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (ch0_yn2_ml_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                         //              (terminated)
		.av_begintransfer         (),                                                                         //              (terminated)
		.av_beginbursttransfer    (),                                                                         //              (terminated)
		.av_burstcount            (),                                                                         //              (terminated)
		.av_byteenable            (),                                                                         //              (terminated)
		.av_readdatavalid         (1'b0),                                                                     //              (terminated)
		.av_waitrequest           (1'b0),                                                                     //              (terminated)
		.av_writebyteenable       (),                                                                         //              (terminated)
		.av_lock                  (),                                                                         //              (terminated)
		.av_clken                 (),                                                                         //              (terminated)
		.uav_clken                (1'b0),                                                                     //              (terminated)
		.av_debugaccess           (),                                                                         //              (terminated)
		.av_outputenable          (),                                                                         //              (terminated)
		.uav_response             (),                                                                         //              (terminated)
		.av_response              (2'b00),                                                                    //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                     //              (terminated)
		.uav_writeresponsevalid   (),                                                                         //              (terminated)
		.av_writeresponserequest  (),                                                                         //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                      //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (22),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ch0_yn2_u_s1_translator (
		.clk                      (clk_clk),                                                                 //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                      //                    reset.reset
		.uav_address              (ch0_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (ch0_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (ch0_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (ch0_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (ch0_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (ch0_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (ch0_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (ch0_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (ch0_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (ch0_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (ch0_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (ch0_yn2_u_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (ch0_yn2_u_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (ch0_yn2_u_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (ch0_yn2_u_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (ch0_yn2_u_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                        //              (terminated)
		.av_begintransfer         (),                                                                        //              (terminated)
		.av_beginbursttransfer    (),                                                                        //              (terminated)
		.av_burstcount            (),                                                                        //              (terminated)
		.av_byteenable            (),                                                                        //              (terminated)
		.av_readdatavalid         (1'b0),                                                                    //              (terminated)
		.av_waitrequest           (1'b0),                                                                    //              (terminated)
		.av_writebyteenable       (),                                                                        //              (terminated)
		.av_lock                  (),                                                                        //              (terminated)
		.av_clken                 (),                                                                        //              (terminated)
		.uav_clken                (1'b0),                                                                    //              (terminated)
		.av_debugaccess           (),                                                                        //              (terminated)
		.av_outputenable          (),                                                                        //              (terminated)
		.uav_response             (),                                                                        //              (terminated)
		.av_response              (2'b00),                                                                   //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                    //              (terminated)
		.uav_writeresponsevalid   (),                                                                        //              (terminated)
		.av_writeresponserequest  (),                                                                        //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                     //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (22),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ch0_yn2_l_s1_translator (
		.clk                      (clk_clk),                                                                 //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                      //                    reset.reset
		.uav_address              (ch0_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (ch0_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (ch0_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (ch0_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (ch0_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (ch0_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (ch0_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (ch0_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (ch0_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (ch0_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (ch0_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (ch0_yn2_l_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (ch0_yn2_l_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (ch0_yn2_l_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (ch0_yn2_l_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (ch0_yn2_l_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                        //              (terminated)
		.av_begintransfer         (),                                                                        //              (terminated)
		.av_beginbursttransfer    (),                                                                        //              (terminated)
		.av_burstcount            (),                                                                        //              (terminated)
		.av_byteenable            (),                                                                        //              (terminated)
		.av_readdatavalid         (1'b0),                                                                    //              (terminated)
		.av_waitrequest           (1'b0),                                                                    //              (terminated)
		.av_writebyteenable       (),                                                                        //              (terminated)
		.av_lock                  (),                                                                        //              (terminated)
		.av_clken                 (),                                                                        //              (terminated)
		.uav_clken                (1'b0),                                                                    //              (terminated)
		.av_debugaccess           (),                                                                        //              (terminated)
		.av_outputenable          (),                                                                        //              (terminated)
		.uav_response             (),                                                                        //              (terminated)
		.av_response              (2'b00),                                                                   //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                    //              (terminated)
		.uav_writeresponsevalid   (),                                                                        //              (terminated)
		.av_writeresponserequest  (),                                                                        //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                     //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (22),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ch0_yn3_l_s1_translator (
		.clk                      (clk_clk),                                                                 //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                      //                    reset.reset
		.uav_address              (ch0_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (ch0_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (ch0_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (ch0_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (ch0_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (ch0_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (ch0_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (ch0_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (ch0_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (ch0_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (ch0_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (ch0_yn3_l_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (ch0_yn3_l_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (ch0_yn3_l_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (ch0_yn3_l_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (ch0_yn3_l_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                        //              (terminated)
		.av_begintransfer         (),                                                                        //              (terminated)
		.av_beginbursttransfer    (),                                                                        //              (terminated)
		.av_burstcount            (),                                                                        //              (terminated)
		.av_byteenable            (),                                                                        //              (terminated)
		.av_readdatavalid         (1'b0),                                                                    //              (terminated)
		.av_waitrequest           (1'b0),                                                                    //              (terminated)
		.av_writebyteenable       (),                                                                        //              (terminated)
		.av_lock                  (),                                                                        //              (terminated)
		.av_clken                 (),                                                                        //              (terminated)
		.uav_clken                (1'b0),                                                                    //              (terminated)
		.av_debugaccess           (),                                                                        //              (terminated)
		.av_outputenable          (),                                                                        //              (terminated)
		.uav_response             (),                                                                        //              (terminated)
		.av_response              (2'b00),                                                                   //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                    //              (terminated)
		.uav_writeresponsevalid   (),                                                                        //              (terminated)
		.av_writeresponserequest  (),                                                                        //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                     //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (22),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ch0_yn3_ml_s1_translator (
		.clk                      (clk_clk),                                                                  //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                       //                    reset.reset
		.uav_address              (ch0_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (ch0_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (ch0_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (ch0_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (ch0_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (ch0_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (ch0_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (ch0_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (ch0_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (ch0_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (ch0_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (ch0_yn3_ml_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (ch0_yn3_ml_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (ch0_yn3_ml_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (ch0_yn3_ml_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (ch0_yn3_ml_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                         //              (terminated)
		.av_begintransfer         (),                                                                         //              (terminated)
		.av_beginbursttransfer    (),                                                                         //              (terminated)
		.av_burstcount            (),                                                                         //              (terminated)
		.av_byteenable            (),                                                                         //              (terminated)
		.av_readdatavalid         (1'b0),                                                                     //              (terminated)
		.av_waitrequest           (1'b0),                                                                     //              (terminated)
		.av_writebyteenable       (),                                                                         //              (terminated)
		.av_lock                  (),                                                                         //              (terminated)
		.av_clken                 (),                                                                         //              (terminated)
		.uav_clken                (1'b0),                                                                     //              (terminated)
		.av_debugaccess           (),                                                                         //              (terminated)
		.av_outputenable          (),                                                                         //              (terminated)
		.uav_response             (),                                                                         //              (terminated)
		.av_response              (2'b00),                                                                    //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                     //              (terminated)
		.uav_writeresponsevalid   (),                                                                         //              (terminated)
		.av_writeresponserequest  (),                                                                         //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                      //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (22),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ch0_yn3_mu_s1_translator (
		.clk                      (clk_clk),                                                                  //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                       //                    reset.reset
		.uav_address              (ch0_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (ch0_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (ch0_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (ch0_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (ch0_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (ch0_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (ch0_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (ch0_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (ch0_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (ch0_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (ch0_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (ch0_yn3_mu_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (ch0_yn3_mu_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (ch0_yn3_mu_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (ch0_yn3_mu_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (ch0_yn3_mu_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                         //              (terminated)
		.av_begintransfer         (),                                                                         //              (terminated)
		.av_beginbursttransfer    (),                                                                         //              (terminated)
		.av_burstcount            (),                                                                         //              (terminated)
		.av_byteenable            (),                                                                         //              (terminated)
		.av_readdatavalid         (1'b0),                                                                     //              (terminated)
		.av_waitrequest           (1'b0),                                                                     //              (terminated)
		.av_writebyteenable       (),                                                                         //              (terminated)
		.av_lock                  (),                                                                         //              (terminated)
		.av_clken                 (),                                                                         //              (terminated)
		.uav_clken                (1'b0),                                                                     //              (terminated)
		.av_debugaccess           (),                                                                         //              (terminated)
		.av_outputenable          (),                                                                         //              (terminated)
		.uav_response             (),                                                                         //              (terminated)
		.av_response              (2'b00),                                                                    //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                     //              (terminated)
		.uav_writeresponsevalid   (),                                                                         //              (terminated)
		.av_writeresponserequest  (),                                                                         //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                      //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (22),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ch0_yn3_u_s1_translator (
		.clk                      (clk_clk),                                                                 //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                      //                    reset.reset
		.uav_address              (ch0_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (ch0_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (ch0_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (ch0_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (ch0_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (ch0_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (ch0_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (ch0_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (ch0_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (ch0_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (ch0_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (ch0_yn3_u_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (ch0_yn3_u_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (ch0_yn3_u_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (ch0_yn3_u_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (ch0_yn3_u_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                        //              (terminated)
		.av_begintransfer         (),                                                                        //              (terminated)
		.av_beginbursttransfer    (),                                                                        //              (terminated)
		.av_burstcount            (),                                                                        //              (terminated)
		.av_byteenable            (),                                                                        //              (terminated)
		.av_readdatavalid         (1'b0),                                                                    //              (terminated)
		.av_waitrequest           (1'b0),                                                                    //              (terminated)
		.av_writebyteenable       (),                                                                        //              (terminated)
		.av_lock                  (),                                                                        //              (terminated)
		.av_clken                 (),                                                                        //              (terminated)
		.uav_clken                (1'b0),                                                                    //              (terminated)
		.av_debugaccess           (),                                                                        //              (terminated)
		.av_outputenable          (),                                                                        //              (terminated)
		.uav_response             (),                                                                        //              (terminated)
		.av_response              (2'b00),                                                                   //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                    //              (terminated)
		.uav_writeresponsevalid   (),                                                                        //              (terminated)
		.av_writeresponserequest  (),                                                                        //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                     //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (22),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ch1_timer_rst_s1_translator (
		.clk                      (clk_clk),                                                                     //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                          //                    reset.reset
		.uav_address              (ch1_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (ch1_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (ch1_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (ch1_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (ch1_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (ch1_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (ch1_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (ch1_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (ch1_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (ch1_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (ch1_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (ch1_timer_rst_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (ch1_timer_rst_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (ch1_timer_rst_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (ch1_timer_rst_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (ch1_timer_rst_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                            //              (terminated)
		.av_begintransfer         (),                                                                            //              (terminated)
		.av_beginbursttransfer    (),                                                                            //              (terminated)
		.av_burstcount            (),                                                                            //              (terminated)
		.av_byteenable            (),                                                                            //              (terminated)
		.av_readdatavalid         (1'b0),                                                                        //              (terminated)
		.av_waitrequest           (1'b0),                                                                        //              (terminated)
		.av_writebyteenable       (),                                                                            //              (terminated)
		.av_lock                  (),                                                                            //              (terminated)
		.av_clken                 (),                                                                            //              (terminated)
		.uav_clken                (1'b0),                                                                        //              (terminated)
		.av_debugaccess           (),                                                                            //              (terminated)
		.av_outputenable          (),                                                                            //              (terminated)
		.uav_response             (),                                                                            //              (terminated)
		.av_response              (2'b00),                                                                       //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                        //              (terminated)
		.uav_writeresponsevalid   (),                                                                            //              (terminated)
		.av_writeresponserequest  (),                                                                            //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                         //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (22),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ch1_thresh_s1_translator (
		.clk                      (clk_clk),                                                                  //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                       //                    reset.reset
		.uav_address              (ch1_thresh_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (ch1_thresh_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (ch1_thresh_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (ch1_thresh_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (ch1_thresh_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (ch1_thresh_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (ch1_thresh_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (ch1_thresh_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (ch1_thresh_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (ch1_thresh_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (ch1_thresh_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (ch1_thresh_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (ch1_thresh_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (ch1_thresh_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (ch1_thresh_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (ch1_thresh_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                         //              (terminated)
		.av_begintransfer         (),                                                                         //              (terminated)
		.av_beginbursttransfer    (),                                                                         //              (terminated)
		.av_burstcount            (),                                                                         //              (terminated)
		.av_byteenable            (),                                                                         //              (terminated)
		.av_readdatavalid         (1'b0),                                                                     //              (terminated)
		.av_waitrequest           (1'b0),                                                                     //              (terminated)
		.av_writebyteenable       (),                                                                         //              (terminated)
		.av_lock                  (),                                                                         //              (terminated)
		.av_clken                 (),                                                                         //              (terminated)
		.uav_clken                (1'b0),                                                                     //              (terminated)
		.av_debugaccess           (),                                                                         //              (terminated)
		.av_outputenable          (),                                                                         //              (terminated)
		.uav_response             (),                                                                         //              (terminated)
		.av_response              (2'b00),                                                                    //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                     //              (terminated)
		.uav_writeresponsevalid   (),                                                                         //              (terminated)
		.av_writeresponserequest  (),                                                                         //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                      //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (22),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ch1_rd_peak_s1_translator (
		.clk                      (clk_clk),                                                                   //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                        //                    reset.reset
		.uav_address              (ch1_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (ch1_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (ch1_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (ch1_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (ch1_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (ch1_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (ch1_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (ch1_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (ch1_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (ch1_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (ch1_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (ch1_rd_peak_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (ch1_rd_peak_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (ch1_rd_peak_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (ch1_rd_peak_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (ch1_rd_peak_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                          //              (terminated)
		.av_begintransfer         (),                                                                          //              (terminated)
		.av_beginbursttransfer    (),                                                                          //              (terminated)
		.av_burstcount            (),                                                                          //              (terminated)
		.av_byteenable            (),                                                                          //              (terminated)
		.av_readdatavalid         (1'b0),                                                                      //              (terminated)
		.av_waitrequest           (1'b0),                                                                      //              (terminated)
		.av_writebyteenable       (),                                                                          //              (terminated)
		.av_lock                  (),                                                                          //              (terminated)
		.av_clken                 (),                                                                          //              (terminated)
		.uav_clken                (1'b0),                                                                      //              (terminated)
		.av_debugaccess           (),                                                                          //              (terminated)
		.av_outputenable          (),                                                                          //              (terminated)
		.uav_response             (),                                                                          //              (terminated)
		.av_response              (2'b00),                                                                     //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                      //              (terminated)
		.uav_writeresponsevalid   (),                                                                          //              (terminated)
		.av_writeresponserequest  (),                                                                          //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                       //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (22),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ch1_peak_found_s1_translator (
		.clk                      (clk_clk),                                                                      //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                           //                    reset.reset
		.uav_address              (ch1_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (ch1_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (ch1_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (ch1_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (ch1_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (ch1_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (ch1_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (ch1_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (ch1_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (ch1_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (ch1_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (ch1_peak_found_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (ch1_peak_found_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (ch1_peak_found_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (ch1_peak_found_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (ch1_peak_found_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                             //              (terminated)
		.av_begintransfer         (),                                                                             //              (terminated)
		.av_beginbursttransfer    (),                                                                             //              (terminated)
		.av_burstcount            (),                                                                             //              (terminated)
		.av_byteenable            (),                                                                             //              (terminated)
		.av_readdatavalid         (1'b0),                                                                         //              (terminated)
		.av_waitrequest           (1'b0),                                                                         //              (terminated)
		.av_writebyteenable       (),                                                                             //              (terminated)
		.av_lock                  (),                                                                             //              (terminated)
		.av_clken                 (),                                                                             //              (terminated)
		.uav_clken                (1'b0),                                                                         //              (terminated)
		.av_debugaccess           (),                                                                             //              (terminated)
		.av_outputenable          (),                                                                             //              (terminated)
		.uav_response             (),                                                                             //              (terminated)
		.av_response              (2'b00),                                                                        //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                         //              (terminated)
		.uav_writeresponsevalid   (),                                                                             //              (terminated)
		.av_writeresponserequest  (),                                                                             //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                          //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (22),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ch1_time_s1_translator (
		.clk                      (clk_clk),                                                                //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                     //                    reset.reset
		.uav_address              (ch1_time_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (ch1_time_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (ch1_time_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (ch1_time_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (ch1_time_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (ch1_time_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (ch1_time_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (ch1_time_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (ch1_time_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (ch1_time_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (ch1_time_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (ch1_time_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (ch1_time_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (ch1_time_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (ch1_time_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (ch1_time_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                       //              (terminated)
		.av_begintransfer         (),                                                                       //              (terminated)
		.av_beginbursttransfer    (),                                                                       //              (terminated)
		.av_burstcount            (),                                                                       //              (terminated)
		.av_byteenable            (),                                                                       //              (terminated)
		.av_readdatavalid         (1'b0),                                                                   //              (terminated)
		.av_waitrequest           (1'b0),                                                                   //              (terminated)
		.av_writebyteenable       (),                                                                       //              (terminated)
		.av_lock                  (),                                                                       //              (terminated)
		.av_clken                 (),                                                                       //              (terminated)
		.uav_clken                (1'b0),                                                                   //              (terminated)
		.av_debugaccess           (),                                                                       //              (terminated)
		.av_outputenable          (),                                                                       //              (terminated)
		.uav_response             (),                                                                       //              (terminated)
		.av_response              (2'b00),                                                                  //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                   //              (terminated)
		.uav_writeresponsevalid   (),                                                                       //              (terminated)
		.av_writeresponserequest  (),                                                                       //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                    //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (22),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ch1_yn1_u_s1_translator (
		.clk                      (clk_clk),                                                                 //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                      //                    reset.reset
		.uav_address              (ch1_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (ch1_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (ch1_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (ch1_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (ch1_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (ch1_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (ch1_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (ch1_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (ch1_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (ch1_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (ch1_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (ch1_yn1_u_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (ch1_yn1_u_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (ch1_yn1_u_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (ch1_yn1_u_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (ch1_yn1_u_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                        //              (terminated)
		.av_begintransfer         (),                                                                        //              (terminated)
		.av_beginbursttransfer    (),                                                                        //              (terminated)
		.av_burstcount            (),                                                                        //              (terminated)
		.av_byteenable            (),                                                                        //              (terminated)
		.av_readdatavalid         (1'b0),                                                                    //              (terminated)
		.av_waitrequest           (1'b0),                                                                    //              (terminated)
		.av_writebyteenable       (),                                                                        //              (terminated)
		.av_lock                  (),                                                                        //              (terminated)
		.av_clken                 (),                                                                        //              (terminated)
		.uav_clken                (1'b0),                                                                    //              (terminated)
		.av_debugaccess           (),                                                                        //              (terminated)
		.av_outputenable          (),                                                                        //              (terminated)
		.uav_response             (),                                                                        //              (terminated)
		.av_response              (2'b00),                                                                   //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                    //              (terminated)
		.uav_writeresponsevalid   (),                                                                        //              (terminated)
		.av_writeresponserequest  (),                                                                        //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                     //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (22),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ch1_yn1_mu_s1_translator (
		.clk                      (clk_clk),                                                                  //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                       //                    reset.reset
		.uav_address              (ch1_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (ch1_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (ch1_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (ch1_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (ch1_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (ch1_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (ch1_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (ch1_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (ch1_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (ch1_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (ch1_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (ch1_yn1_mu_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (ch1_yn1_mu_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (ch1_yn1_mu_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (ch1_yn1_mu_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (ch1_yn1_mu_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                         //              (terminated)
		.av_begintransfer         (),                                                                         //              (terminated)
		.av_beginbursttransfer    (),                                                                         //              (terminated)
		.av_burstcount            (),                                                                         //              (terminated)
		.av_byteenable            (),                                                                         //              (terminated)
		.av_readdatavalid         (1'b0),                                                                     //              (terminated)
		.av_waitrequest           (1'b0),                                                                     //              (terminated)
		.av_writebyteenable       (),                                                                         //              (terminated)
		.av_lock                  (),                                                                         //              (terminated)
		.av_clken                 (),                                                                         //              (terminated)
		.uav_clken                (1'b0),                                                                     //              (terminated)
		.av_debugaccess           (),                                                                         //              (terminated)
		.av_outputenable          (),                                                                         //              (terminated)
		.uav_response             (),                                                                         //              (terminated)
		.av_response              (2'b00),                                                                    //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                     //              (terminated)
		.uav_writeresponsevalid   (),                                                                         //              (terminated)
		.av_writeresponserequest  (),                                                                         //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                      //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (22),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ch1_yn1_ml_s1_translator (
		.clk                      (clk_clk),                                                                  //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                       //                    reset.reset
		.uav_address              (ch1_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (ch1_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (ch1_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (ch1_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (ch1_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (ch1_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (ch1_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (ch1_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (ch1_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (ch1_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (ch1_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (ch1_yn1_ml_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (ch1_yn1_ml_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (ch1_yn1_ml_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (ch1_yn1_ml_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (ch1_yn1_ml_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                         //              (terminated)
		.av_begintransfer         (),                                                                         //              (terminated)
		.av_beginbursttransfer    (),                                                                         //              (terminated)
		.av_burstcount            (),                                                                         //              (terminated)
		.av_byteenable            (),                                                                         //              (terminated)
		.av_readdatavalid         (1'b0),                                                                     //              (terminated)
		.av_waitrequest           (1'b0),                                                                     //              (terminated)
		.av_writebyteenable       (),                                                                         //              (terminated)
		.av_lock                  (),                                                                         //              (terminated)
		.av_clken                 (),                                                                         //              (terminated)
		.uav_clken                (1'b0),                                                                     //              (terminated)
		.av_debugaccess           (),                                                                         //              (terminated)
		.av_outputenable          (),                                                                         //              (terminated)
		.uav_response             (),                                                                         //              (terminated)
		.av_response              (2'b00),                                                                    //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                     //              (terminated)
		.uav_writeresponsevalid   (),                                                                         //              (terminated)
		.av_writeresponserequest  (),                                                                         //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                      //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (22),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ch1_yn1_l_s1_translator (
		.clk                      (clk_clk),                                                                 //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                      //                    reset.reset
		.uav_address              (ch1_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (ch1_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (ch1_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (ch1_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (ch1_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (ch1_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (ch1_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (ch1_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (ch1_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (ch1_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (ch1_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (ch1_yn1_l_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (ch1_yn1_l_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (ch1_yn1_l_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (ch1_yn1_l_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (ch1_yn1_l_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                        //              (terminated)
		.av_begintransfer         (),                                                                        //              (terminated)
		.av_beginbursttransfer    (),                                                                        //              (terminated)
		.av_burstcount            (),                                                                        //              (terminated)
		.av_byteenable            (),                                                                        //              (terminated)
		.av_readdatavalid         (1'b0),                                                                    //              (terminated)
		.av_waitrequest           (1'b0),                                                                    //              (terminated)
		.av_writebyteenable       (),                                                                        //              (terminated)
		.av_lock                  (),                                                                        //              (terminated)
		.av_clken                 (),                                                                        //              (terminated)
		.uav_clken                (1'b0),                                                                    //              (terminated)
		.av_debugaccess           (),                                                                        //              (terminated)
		.av_outputenable          (),                                                                        //              (terminated)
		.uav_response             (),                                                                        //              (terminated)
		.av_response              (2'b00),                                                                   //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                    //              (terminated)
		.uav_writeresponsevalid   (),                                                                        //              (terminated)
		.av_writeresponserequest  (),                                                                        //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                     //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (22),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ch1_yn2_u_s1_translator (
		.clk                      (clk_clk),                                                                 //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                      //                    reset.reset
		.uav_address              (ch1_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (ch1_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (ch1_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (ch1_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (ch1_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (ch1_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (ch1_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (ch1_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (ch1_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (ch1_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (ch1_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (ch1_yn2_u_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (ch1_yn2_u_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (ch1_yn2_u_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (ch1_yn2_u_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (ch1_yn2_u_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                        //              (terminated)
		.av_begintransfer         (),                                                                        //              (terminated)
		.av_beginbursttransfer    (),                                                                        //              (terminated)
		.av_burstcount            (),                                                                        //              (terminated)
		.av_byteenable            (),                                                                        //              (terminated)
		.av_readdatavalid         (1'b0),                                                                    //              (terminated)
		.av_waitrequest           (1'b0),                                                                    //              (terminated)
		.av_writebyteenable       (),                                                                        //              (terminated)
		.av_lock                  (),                                                                        //              (terminated)
		.av_clken                 (),                                                                        //              (terminated)
		.uav_clken                (1'b0),                                                                    //              (terminated)
		.av_debugaccess           (),                                                                        //              (terminated)
		.av_outputenable          (),                                                                        //              (terminated)
		.uav_response             (),                                                                        //              (terminated)
		.av_response              (2'b00),                                                                   //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                    //              (terminated)
		.uav_writeresponsevalid   (),                                                                        //              (terminated)
		.av_writeresponserequest  (),                                                                        //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                     //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (22),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ch1_yn2_mu_s1_translator (
		.clk                      (clk_clk),                                                                  //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                       //                    reset.reset
		.uav_address              (ch1_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (ch1_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (ch1_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (ch1_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (ch1_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (ch1_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (ch1_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (ch1_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (ch1_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (ch1_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (ch1_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (ch1_yn2_mu_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (ch1_yn2_mu_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (ch1_yn2_mu_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (ch1_yn2_mu_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (ch1_yn2_mu_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                         //              (terminated)
		.av_begintransfer         (),                                                                         //              (terminated)
		.av_beginbursttransfer    (),                                                                         //              (terminated)
		.av_burstcount            (),                                                                         //              (terminated)
		.av_byteenable            (),                                                                         //              (terminated)
		.av_readdatavalid         (1'b0),                                                                     //              (terminated)
		.av_waitrequest           (1'b0),                                                                     //              (terminated)
		.av_writebyteenable       (),                                                                         //              (terminated)
		.av_lock                  (),                                                                         //              (terminated)
		.av_clken                 (),                                                                         //              (terminated)
		.uav_clken                (1'b0),                                                                     //              (terminated)
		.av_debugaccess           (),                                                                         //              (terminated)
		.av_outputenable          (),                                                                         //              (terminated)
		.uav_response             (),                                                                         //              (terminated)
		.av_response              (2'b00),                                                                    //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                     //              (terminated)
		.uav_writeresponsevalid   (),                                                                         //              (terminated)
		.av_writeresponserequest  (),                                                                         //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                      //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (22),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ch1_yn2_ml_s1_translator (
		.clk                      (clk_clk),                                                                  //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                       //                    reset.reset
		.uav_address              (ch1_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (ch1_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (ch1_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (ch1_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (ch1_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (ch1_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (ch1_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (ch1_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (ch1_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (ch1_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (ch1_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (ch1_yn2_ml_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (ch1_yn2_ml_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (ch1_yn2_ml_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (ch1_yn2_ml_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (ch1_yn2_ml_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                         //              (terminated)
		.av_begintransfer         (),                                                                         //              (terminated)
		.av_beginbursttransfer    (),                                                                         //              (terminated)
		.av_burstcount            (),                                                                         //              (terminated)
		.av_byteenable            (),                                                                         //              (terminated)
		.av_readdatavalid         (1'b0),                                                                     //              (terminated)
		.av_waitrequest           (1'b0),                                                                     //              (terminated)
		.av_writebyteenable       (),                                                                         //              (terminated)
		.av_lock                  (),                                                                         //              (terminated)
		.av_clken                 (),                                                                         //              (terminated)
		.uav_clken                (1'b0),                                                                     //              (terminated)
		.av_debugaccess           (),                                                                         //              (terminated)
		.av_outputenable          (),                                                                         //              (terminated)
		.uav_response             (),                                                                         //              (terminated)
		.av_response              (2'b00),                                                                    //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                     //              (terminated)
		.uav_writeresponsevalid   (),                                                                         //              (terminated)
		.av_writeresponserequest  (),                                                                         //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                      //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (22),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ch1_yn2_l_s1_translator (
		.clk                      (clk_clk),                                                                 //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                      //                    reset.reset
		.uav_address              (ch1_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (ch1_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (ch1_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (ch1_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (ch1_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (ch1_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (ch1_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (ch1_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (ch1_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (ch1_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (ch1_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (ch1_yn2_l_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (ch1_yn2_l_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (ch1_yn2_l_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (ch1_yn2_l_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (ch1_yn2_l_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                        //              (terminated)
		.av_begintransfer         (),                                                                        //              (terminated)
		.av_beginbursttransfer    (),                                                                        //              (terminated)
		.av_burstcount            (),                                                                        //              (terminated)
		.av_byteenable            (),                                                                        //              (terminated)
		.av_readdatavalid         (1'b0),                                                                    //              (terminated)
		.av_waitrequest           (1'b0),                                                                    //              (terminated)
		.av_writebyteenable       (),                                                                        //              (terminated)
		.av_lock                  (),                                                                        //              (terminated)
		.av_clken                 (),                                                                        //              (terminated)
		.uav_clken                (1'b0),                                                                    //              (terminated)
		.av_debugaccess           (),                                                                        //              (terminated)
		.av_outputenable          (),                                                                        //              (terminated)
		.uav_response             (),                                                                        //              (terminated)
		.av_response              (2'b00),                                                                   //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                    //              (terminated)
		.uav_writeresponsevalid   (),                                                                        //              (terminated)
		.av_writeresponserequest  (),                                                                        //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                     //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (22),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ch1_yn3_u_s1_translator (
		.clk                      (clk_clk),                                                                 //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                      //                    reset.reset
		.uav_address              (ch1_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (ch1_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (ch1_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (ch1_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (ch1_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (ch1_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (ch1_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (ch1_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (ch1_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (ch1_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (ch1_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (ch1_yn3_u_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (ch1_yn3_u_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (ch1_yn3_u_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (ch1_yn3_u_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (ch1_yn3_u_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                        //              (terminated)
		.av_begintransfer         (),                                                                        //              (terminated)
		.av_beginbursttransfer    (),                                                                        //              (terminated)
		.av_burstcount            (),                                                                        //              (terminated)
		.av_byteenable            (),                                                                        //              (terminated)
		.av_readdatavalid         (1'b0),                                                                    //              (terminated)
		.av_waitrequest           (1'b0),                                                                    //              (terminated)
		.av_writebyteenable       (),                                                                        //              (terminated)
		.av_lock                  (),                                                                        //              (terminated)
		.av_clken                 (),                                                                        //              (terminated)
		.uav_clken                (1'b0),                                                                    //              (terminated)
		.av_debugaccess           (),                                                                        //              (terminated)
		.av_outputenable          (),                                                                        //              (terminated)
		.uav_response             (),                                                                        //              (terminated)
		.av_response              (2'b00),                                                                   //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                    //              (terminated)
		.uav_writeresponsevalid   (),                                                                        //              (terminated)
		.av_writeresponserequest  (),                                                                        //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                     //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (22),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ch1_yn3_mu_s1_translator (
		.clk                      (clk_clk),                                                                  //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                       //                    reset.reset
		.uav_address              (ch1_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (ch1_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (ch1_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (ch1_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (ch1_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (ch1_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (ch1_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (ch1_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (ch1_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (ch1_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (ch1_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (ch1_yn3_mu_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (ch1_yn3_mu_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (ch1_yn3_mu_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (ch1_yn3_mu_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (ch1_yn3_mu_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                         //              (terminated)
		.av_begintransfer         (),                                                                         //              (terminated)
		.av_beginbursttransfer    (),                                                                         //              (terminated)
		.av_burstcount            (),                                                                         //              (terminated)
		.av_byteenable            (),                                                                         //              (terminated)
		.av_readdatavalid         (1'b0),                                                                     //              (terminated)
		.av_waitrequest           (1'b0),                                                                     //              (terminated)
		.av_writebyteenable       (),                                                                         //              (terminated)
		.av_lock                  (),                                                                         //              (terminated)
		.av_clken                 (),                                                                         //              (terminated)
		.uav_clken                (1'b0),                                                                     //              (terminated)
		.av_debugaccess           (),                                                                         //              (terminated)
		.av_outputenable          (),                                                                         //              (terminated)
		.uav_response             (),                                                                         //              (terminated)
		.av_response              (2'b00),                                                                    //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                     //              (terminated)
		.uav_writeresponsevalid   (),                                                                         //              (terminated)
		.av_writeresponserequest  (),                                                                         //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                      //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (22),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ch1_yn3_ml_s1_translator (
		.clk                      (clk_clk),                                                                  //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                       //                    reset.reset
		.uav_address              (ch1_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (ch1_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (ch1_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (ch1_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (ch1_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (ch1_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (ch1_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (ch1_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (ch1_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (ch1_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (ch1_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (ch1_yn3_ml_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (ch1_yn3_ml_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (ch1_yn3_ml_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (ch1_yn3_ml_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (ch1_yn3_ml_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                         //              (terminated)
		.av_begintransfer         (),                                                                         //              (terminated)
		.av_beginbursttransfer    (),                                                                         //              (terminated)
		.av_burstcount            (),                                                                         //              (terminated)
		.av_byteenable            (),                                                                         //              (terminated)
		.av_readdatavalid         (1'b0),                                                                     //              (terminated)
		.av_waitrequest           (1'b0),                                                                     //              (terminated)
		.av_writebyteenable       (),                                                                         //              (terminated)
		.av_lock                  (),                                                                         //              (terminated)
		.av_clken                 (),                                                                         //              (terminated)
		.uav_clken                (1'b0),                                                                     //              (terminated)
		.av_debugaccess           (),                                                                         //              (terminated)
		.av_outputenable          (),                                                                         //              (terminated)
		.uav_response             (),                                                                         //              (terminated)
		.av_response              (2'b00),                                                                    //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                     //              (terminated)
		.uav_writeresponsevalid   (),                                                                         //              (terminated)
		.av_writeresponserequest  (),                                                                         //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                      //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (22),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ch1_yn3_l_s1_translator (
		.clk                      (clk_clk),                                                                 //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                      //                    reset.reset
		.uav_address              (ch1_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (ch1_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (ch1_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (ch1_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (ch1_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (ch1_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (ch1_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (ch1_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (ch1_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (ch1_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (ch1_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (ch1_yn3_l_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (ch1_yn3_l_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (ch1_yn3_l_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (ch1_yn3_l_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (ch1_yn3_l_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                        //              (terminated)
		.av_begintransfer         (),                                                                        //              (terminated)
		.av_beginbursttransfer    (),                                                                        //              (terminated)
		.av_burstcount            (),                                                                        //              (terminated)
		.av_byteenable            (),                                                                        //              (terminated)
		.av_readdatavalid         (1'b0),                                                                    //              (terminated)
		.av_waitrequest           (1'b0),                                                                    //              (terminated)
		.av_writebyteenable       (),                                                                        //              (terminated)
		.av_lock                  (),                                                                        //              (terminated)
		.av_clken                 (),                                                                        //              (terminated)
		.uav_clken                (1'b0),                                                                    //              (terminated)
		.av_debugaccess           (),                                                                        //              (terminated)
		.av_outputenable          (),                                                                        //              (terminated)
		.uav_response             (),                                                                        //              (terminated)
		.av_response              (2'b00),                                                                   //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                    //              (terminated)
		.uav_writeresponsevalid   (),                                                                        //              (terminated)
		.av_writeresponserequest  (),                                                                        //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                     //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (22),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ch2_timer_rst_s1_translator (
		.clk                      (clk_clk),                                                                     //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                          //                    reset.reset
		.uav_address              (ch2_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (ch2_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (ch2_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (ch2_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (ch2_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (ch2_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (ch2_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (ch2_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (ch2_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (ch2_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (ch2_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (ch2_timer_rst_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (ch2_timer_rst_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (ch2_timer_rst_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (ch2_timer_rst_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (ch2_timer_rst_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                            //              (terminated)
		.av_begintransfer         (),                                                                            //              (terminated)
		.av_beginbursttransfer    (),                                                                            //              (terminated)
		.av_burstcount            (),                                                                            //              (terminated)
		.av_byteenable            (),                                                                            //              (terminated)
		.av_readdatavalid         (1'b0),                                                                        //              (terminated)
		.av_waitrequest           (1'b0),                                                                        //              (terminated)
		.av_writebyteenable       (),                                                                            //              (terminated)
		.av_lock                  (),                                                                            //              (terminated)
		.av_clken                 (),                                                                            //              (terminated)
		.uav_clken                (1'b0),                                                                        //              (terminated)
		.av_debugaccess           (),                                                                            //              (terminated)
		.av_outputenable          (),                                                                            //              (terminated)
		.uav_response             (),                                                                            //              (terminated)
		.av_response              (2'b00),                                                                       //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                        //              (terminated)
		.uav_writeresponsevalid   (),                                                                            //              (terminated)
		.av_writeresponserequest  (),                                                                            //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                         //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (22),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ch2_thresh_s1_translator (
		.clk                      (clk_clk),                                                                  //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                       //                    reset.reset
		.uav_address              (ch2_thresh_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (ch2_thresh_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (ch2_thresh_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (ch2_thresh_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (ch2_thresh_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (ch2_thresh_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (ch2_thresh_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (ch2_thresh_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (ch2_thresh_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (ch2_thresh_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (ch2_thresh_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (ch2_thresh_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (ch2_thresh_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (ch2_thresh_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (ch2_thresh_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (ch2_thresh_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                         //              (terminated)
		.av_begintransfer         (),                                                                         //              (terminated)
		.av_beginbursttransfer    (),                                                                         //              (terminated)
		.av_burstcount            (),                                                                         //              (terminated)
		.av_byteenable            (),                                                                         //              (terminated)
		.av_readdatavalid         (1'b0),                                                                     //              (terminated)
		.av_waitrequest           (1'b0),                                                                     //              (terminated)
		.av_writebyteenable       (),                                                                         //              (terminated)
		.av_lock                  (),                                                                         //              (terminated)
		.av_clken                 (),                                                                         //              (terminated)
		.uav_clken                (1'b0),                                                                     //              (terminated)
		.av_debugaccess           (),                                                                         //              (terminated)
		.av_outputenable          (),                                                                         //              (terminated)
		.uav_response             (),                                                                         //              (terminated)
		.av_response              (2'b00),                                                                    //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                     //              (terminated)
		.uav_writeresponsevalid   (),                                                                         //              (terminated)
		.av_writeresponserequest  (),                                                                         //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                      //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (22),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ch2_rd_peak_s1_translator (
		.clk                      (clk_clk),                                                                   //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                        //                    reset.reset
		.uav_address              (ch2_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (ch2_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (ch2_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (ch2_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (ch2_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (ch2_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (ch2_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (ch2_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (ch2_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (ch2_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (ch2_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (ch2_rd_peak_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (ch2_rd_peak_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (ch2_rd_peak_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (ch2_rd_peak_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (ch2_rd_peak_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                          //              (terminated)
		.av_begintransfer         (),                                                                          //              (terminated)
		.av_beginbursttransfer    (),                                                                          //              (terminated)
		.av_burstcount            (),                                                                          //              (terminated)
		.av_byteenable            (),                                                                          //              (terminated)
		.av_readdatavalid         (1'b0),                                                                      //              (terminated)
		.av_waitrequest           (1'b0),                                                                      //              (terminated)
		.av_writebyteenable       (),                                                                          //              (terminated)
		.av_lock                  (),                                                                          //              (terminated)
		.av_clken                 (),                                                                          //              (terminated)
		.uav_clken                (1'b0),                                                                      //              (terminated)
		.av_debugaccess           (),                                                                          //              (terminated)
		.av_outputenable          (),                                                                          //              (terminated)
		.uav_response             (),                                                                          //              (terminated)
		.av_response              (2'b00),                                                                     //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                      //              (terminated)
		.uav_writeresponsevalid   (),                                                                          //              (terminated)
		.av_writeresponserequest  (),                                                                          //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                       //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (22),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ch2_peak_found_s1_translator (
		.clk                      (clk_clk),                                                                      //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                           //                    reset.reset
		.uav_address              (ch2_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (ch2_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (ch2_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (ch2_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (ch2_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (ch2_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (ch2_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (ch2_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (ch2_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (ch2_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (ch2_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (ch2_peak_found_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (ch2_peak_found_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (ch2_peak_found_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (ch2_peak_found_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (ch2_peak_found_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                             //              (terminated)
		.av_begintransfer         (),                                                                             //              (terminated)
		.av_beginbursttransfer    (),                                                                             //              (terminated)
		.av_burstcount            (),                                                                             //              (terminated)
		.av_byteenable            (),                                                                             //              (terminated)
		.av_readdatavalid         (1'b0),                                                                         //              (terminated)
		.av_waitrequest           (1'b0),                                                                         //              (terminated)
		.av_writebyteenable       (),                                                                             //              (terminated)
		.av_lock                  (),                                                                             //              (terminated)
		.av_clken                 (),                                                                             //              (terminated)
		.uav_clken                (1'b0),                                                                         //              (terminated)
		.av_debugaccess           (),                                                                             //              (terminated)
		.av_outputenable          (),                                                                             //              (terminated)
		.uav_response             (),                                                                             //              (terminated)
		.av_response              (2'b00),                                                                        //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                         //              (terminated)
		.uav_writeresponsevalid   (),                                                                             //              (terminated)
		.av_writeresponserequest  (),                                                                             //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                          //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (22),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ch2_time_s1_translator (
		.clk                      (clk_clk),                                                                //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                     //                    reset.reset
		.uav_address              (ch2_time_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (ch2_time_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (ch2_time_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (ch2_time_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (ch2_time_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (ch2_time_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (ch2_time_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (ch2_time_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (ch2_time_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (ch2_time_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (ch2_time_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (ch2_time_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (ch2_time_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (ch2_time_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (ch2_time_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (ch2_time_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                       //              (terminated)
		.av_begintransfer         (),                                                                       //              (terminated)
		.av_beginbursttransfer    (),                                                                       //              (terminated)
		.av_burstcount            (),                                                                       //              (terminated)
		.av_byteenable            (),                                                                       //              (terminated)
		.av_readdatavalid         (1'b0),                                                                   //              (terminated)
		.av_waitrequest           (1'b0),                                                                   //              (terminated)
		.av_writebyteenable       (),                                                                       //              (terminated)
		.av_lock                  (),                                                                       //              (terminated)
		.av_clken                 (),                                                                       //              (terminated)
		.uav_clken                (1'b0),                                                                   //              (terminated)
		.av_debugaccess           (),                                                                       //              (terminated)
		.av_outputenable          (),                                                                       //              (terminated)
		.uav_response             (),                                                                       //              (terminated)
		.av_response              (2'b00),                                                                  //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                   //              (terminated)
		.uav_writeresponsevalid   (),                                                                       //              (terminated)
		.av_writeresponserequest  (),                                                                       //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                    //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (22),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ch2_yn1_u_s1_translator (
		.clk                      (clk_clk),                                                                 //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                      //                    reset.reset
		.uav_address              (ch2_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (ch2_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (ch2_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (ch2_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (ch2_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (ch2_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (ch2_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (ch2_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (ch2_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (ch2_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (ch2_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (ch2_yn1_u_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (ch2_yn1_u_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (ch2_yn1_u_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (ch2_yn1_u_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (ch2_yn1_u_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                        //              (terminated)
		.av_begintransfer         (),                                                                        //              (terminated)
		.av_beginbursttransfer    (),                                                                        //              (terminated)
		.av_burstcount            (),                                                                        //              (terminated)
		.av_byteenable            (),                                                                        //              (terminated)
		.av_readdatavalid         (1'b0),                                                                    //              (terminated)
		.av_waitrequest           (1'b0),                                                                    //              (terminated)
		.av_writebyteenable       (),                                                                        //              (terminated)
		.av_lock                  (),                                                                        //              (terminated)
		.av_clken                 (),                                                                        //              (terminated)
		.uav_clken                (1'b0),                                                                    //              (terminated)
		.av_debugaccess           (),                                                                        //              (terminated)
		.av_outputenable          (),                                                                        //              (terminated)
		.uav_response             (),                                                                        //              (terminated)
		.av_response              (2'b00),                                                                   //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                    //              (terminated)
		.uav_writeresponsevalid   (),                                                                        //              (terminated)
		.av_writeresponserequest  (),                                                                        //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                     //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (22),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ch2_yn1_mu_s1_translator (
		.clk                      (clk_clk),                                                                  //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                       //                    reset.reset
		.uav_address              (ch2_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (ch2_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (ch2_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (ch2_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (ch2_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (ch2_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (ch2_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (ch2_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (ch2_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (ch2_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (ch2_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (ch2_yn1_mu_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (ch2_yn1_mu_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (ch2_yn1_mu_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (ch2_yn1_mu_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (ch2_yn1_mu_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                         //              (terminated)
		.av_begintransfer         (),                                                                         //              (terminated)
		.av_beginbursttransfer    (),                                                                         //              (terminated)
		.av_burstcount            (),                                                                         //              (terminated)
		.av_byteenable            (),                                                                         //              (terminated)
		.av_readdatavalid         (1'b0),                                                                     //              (terminated)
		.av_waitrequest           (1'b0),                                                                     //              (terminated)
		.av_writebyteenable       (),                                                                         //              (terminated)
		.av_lock                  (),                                                                         //              (terminated)
		.av_clken                 (),                                                                         //              (terminated)
		.uav_clken                (1'b0),                                                                     //              (terminated)
		.av_debugaccess           (),                                                                         //              (terminated)
		.av_outputenable          (),                                                                         //              (terminated)
		.uav_response             (),                                                                         //              (terminated)
		.av_response              (2'b00),                                                                    //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                     //              (terminated)
		.uav_writeresponsevalid   (),                                                                         //              (terminated)
		.av_writeresponserequest  (),                                                                         //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                      //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (22),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ch2_yn1_ml_s1_translator (
		.clk                      (clk_clk),                                                                  //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                       //                    reset.reset
		.uav_address              (ch2_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (ch2_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (ch2_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (ch2_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (ch2_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (ch2_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (ch2_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (ch2_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (ch2_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (ch2_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (ch2_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (ch2_yn1_ml_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (ch2_yn1_ml_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (ch2_yn1_ml_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (ch2_yn1_ml_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (ch2_yn1_ml_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                         //              (terminated)
		.av_begintransfer         (),                                                                         //              (terminated)
		.av_beginbursttransfer    (),                                                                         //              (terminated)
		.av_burstcount            (),                                                                         //              (terminated)
		.av_byteenable            (),                                                                         //              (terminated)
		.av_readdatavalid         (1'b0),                                                                     //              (terminated)
		.av_waitrequest           (1'b0),                                                                     //              (terminated)
		.av_writebyteenable       (),                                                                         //              (terminated)
		.av_lock                  (),                                                                         //              (terminated)
		.av_clken                 (),                                                                         //              (terminated)
		.uav_clken                (1'b0),                                                                     //              (terminated)
		.av_debugaccess           (),                                                                         //              (terminated)
		.av_outputenable          (),                                                                         //              (terminated)
		.uav_response             (),                                                                         //              (terminated)
		.av_response              (2'b00),                                                                    //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                     //              (terminated)
		.uav_writeresponsevalid   (),                                                                         //              (terminated)
		.av_writeresponserequest  (),                                                                         //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                      //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (22),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ch2_yn1_l_s1_translator (
		.clk                      (clk_clk),                                                                 //                      clk.clk
		.reset                    (nios_cpu_jtag_debug_module_reset_reset),                                  //                    reset.reset
		.uav_address              (ch2_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (ch2_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (ch2_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (ch2_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (ch2_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (ch2_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (ch2_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (ch2_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (ch2_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (ch2_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (ch2_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (ch2_yn1_l_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (ch2_yn1_l_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (ch2_yn1_l_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (ch2_yn1_l_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (ch2_yn1_l_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                        //              (terminated)
		.av_begintransfer         (),                                                                        //              (terminated)
		.av_beginbursttransfer    (),                                                                        //              (terminated)
		.av_burstcount            (),                                                                        //              (terminated)
		.av_byteenable            (),                                                                        //              (terminated)
		.av_readdatavalid         (1'b0),                                                                    //              (terminated)
		.av_waitrequest           (1'b0),                                                                    //              (terminated)
		.av_writebyteenable       (),                                                                        //              (terminated)
		.av_lock                  (),                                                                        //              (terminated)
		.av_clken                 (),                                                                        //              (terminated)
		.uav_clken                (1'b0),                                                                    //              (terminated)
		.av_debugaccess           (),                                                                        //              (terminated)
		.av_outputenable          (),                                                                        //              (terminated)
		.uav_response             (),                                                                        //              (terminated)
		.av_response              (2'b00),                                                                   //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                    //              (terminated)
		.uav_writeresponsevalid   (),                                                                        //              (terminated)
		.av_writeresponserequest  (),                                                                        //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                     //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (22),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ch2_yn2_u_s1_translator (
		.clk                      (clk_clk),                                                                 //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                      //                    reset.reset
		.uav_address              (ch2_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (ch2_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (ch2_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (ch2_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (ch2_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (ch2_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (ch2_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (ch2_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (ch2_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (ch2_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (ch2_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (ch2_yn2_u_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (ch2_yn2_u_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (ch2_yn2_u_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (ch2_yn2_u_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (ch2_yn2_u_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                        //              (terminated)
		.av_begintransfer         (),                                                                        //              (terminated)
		.av_beginbursttransfer    (),                                                                        //              (terminated)
		.av_burstcount            (),                                                                        //              (terminated)
		.av_byteenable            (),                                                                        //              (terminated)
		.av_readdatavalid         (1'b0),                                                                    //              (terminated)
		.av_waitrequest           (1'b0),                                                                    //              (terminated)
		.av_writebyteenable       (),                                                                        //              (terminated)
		.av_lock                  (),                                                                        //              (terminated)
		.av_clken                 (),                                                                        //              (terminated)
		.uav_clken                (1'b0),                                                                    //              (terminated)
		.av_debugaccess           (),                                                                        //              (terminated)
		.av_outputenable          (),                                                                        //              (terminated)
		.uav_response             (),                                                                        //              (terminated)
		.av_response              (2'b00),                                                                   //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                    //              (terminated)
		.uav_writeresponsevalid   (),                                                                        //              (terminated)
		.av_writeresponserequest  (),                                                                        //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                     //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (22),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ch2_yn2_mu_s1_translator (
		.clk                      (clk_clk),                                                                  //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                       //                    reset.reset
		.uav_address              (ch2_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (ch2_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (ch2_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (ch2_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (ch2_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (ch2_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (ch2_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (ch2_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (ch2_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (ch2_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (ch2_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (ch2_yn2_mu_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (ch2_yn2_mu_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (ch2_yn2_mu_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (ch2_yn2_mu_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (ch2_yn2_mu_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                         //              (terminated)
		.av_begintransfer         (),                                                                         //              (terminated)
		.av_beginbursttransfer    (),                                                                         //              (terminated)
		.av_burstcount            (),                                                                         //              (terminated)
		.av_byteenable            (),                                                                         //              (terminated)
		.av_readdatavalid         (1'b0),                                                                     //              (terminated)
		.av_waitrequest           (1'b0),                                                                     //              (terminated)
		.av_writebyteenable       (),                                                                         //              (terminated)
		.av_lock                  (),                                                                         //              (terminated)
		.av_clken                 (),                                                                         //              (terminated)
		.uav_clken                (1'b0),                                                                     //              (terminated)
		.av_debugaccess           (),                                                                         //              (terminated)
		.av_outputenable          (),                                                                         //              (terminated)
		.uav_response             (),                                                                         //              (terminated)
		.av_response              (2'b00),                                                                    //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                     //              (terminated)
		.uav_writeresponsevalid   (),                                                                         //              (terminated)
		.av_writeresponserequest  (),                                                                         //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                      //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (22),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ch2_yn2_ml_s1_translator (
		.clk                      (clk_clk),                                                                  //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                       //                    reset.reset
		.uav_address              (ch2_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (ch2_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (ch2_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (ch2_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (ch2_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (ch2_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (ch2_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (ch2_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (ch2_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (ch2_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (ch2_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (ch2_yn2_ml_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (ch2_yn2_ml_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (ch2_yn2_ml_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (ch2_yn2_ml_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (ch2_yn2_ml_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                         //              (terminated)
		.av_begintransfer         (),                                                                         //              (terminated)
		.av_beginbursttransfer    (),                                                                         //              (terminated)
		.av_burstcount            (),                                                                         //              (terminated)
		.av_byteenable            (),                                                                         //              (terminated)
		.av_readdatavalid         (1'b0),                                                                     //              (terminated)
		.av_waitrequest           (1'b0),                                                                     //              (terminated)
		.av_writebyteenable       (),                                                                         //              (terminated)
		.av_lock                  (),                                                                         //              (terminated)
		.av_clken                 (),                                                                         //              (terminated)
		.uav_clken                (1'b0),                                                                     //              (terminated)
		.av_debugaccess           (),                                                                         //              (terminated)
		.av_outputenable          (),                                                                         //              (terminated)
		.uav_response             (),                                                                         //              (terminated)
		.av_response              (2'b00),                                                                    //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                     //              (terminated)
		.uav_writeresponsevalid   (),                                                                         //              (terminated)
		.av_writeresponserequest  (),                                                                         //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                      //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (22),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ch2_yn2_l_s1_translator (
		.clk                      (clk_clk),                                                                 //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                      //                    reset.reset
		.uav_address              (ch2_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (ch2_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (ch2_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (ch2_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (ch2_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (ch2_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (ch2_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (ch2_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (ch2_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (ch2_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (ch2_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (ch2_yn2_l_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (ch2_yn2_l_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (ch2_yn2_l_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (ch2_yn2_l_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (ch2_yn2_l_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                        //              (terminated)
		.av_begintransfer         (),                                                                        //              (terminated)
		.av_beginbursttransfer    (),                                                                        //              (terminated)
		.av_burstcount            (),                                                                        //              (terminated)
		.av_byteenable            (),                                                                        //              (terminated)
		.av_readdatavalid         (1'b0),                                                                    //              (terminated)
		.av_waitrequest           (1'b0),                                                                    //              (terminated)
		.av_writebyteenable       (),                                                                        //              (terminated)
		.av_lock                  (),                                                                        //              (terminated)
		.av_clken                 (),                                                                        //              (terminated)
		.uav_clken                (1'b0),                                                                    //              (terminated)
		.av_debugaccess           (),                                                                        //              (terminated)
		.av_outputenable          (),                                                                        //              (terminated)
		.uav_response             (),                                                                        //              (terminated)
		.av_response              (2'b00),                                                                   //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                    //              (terminated)
		.uav_writeresponsevalid   (),                                                                        //              (terminated)
		.av_writeresponserequest  (),                                                                        //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                     //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (22),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ch2_yn3_u_s1_translator (
		.clk                      (clk_clk),                                                                 //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                      //                    reset.reset
		.uav_address              (ch2_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (ch2_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (ch2_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (ch2_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (ch2_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (ch2_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (ch2_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (ch2_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (ch2_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (ch2_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (ch2_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (ch2_yn3_u_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (ch2_yn3_u_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (ch2_yn3_u_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (ch2_yn3_u_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (ch2_yn3_u_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                        //              (terminated)
		.av_begintransfer         (),                                                                        //              (terminated)
		.av_beginbursttransfer    (),                                                                        //              (terminated)
		.av_burstcount            (),                                                                        //              (terminated)
		.av_byteenable            (),                                                                        //              (terminated)
		.av_readdatavalid         (1'b0),                                                                    //              (terminated)
		.av_waitrequest           (1'b0),                                                                    //              (terminated)
		.av_writebyteenable       (),                                                                        //              (terminated)
		.av_lock                  (),                                                                        //              (terminated)
		.av_clken                 (),                                                                        //              (terminated)
		.uav_clken                (1'b0),                                                                    //              (terminated)
		.av_debugaccess           (),                                                                        //              (terminated)
		.av_outputenable          (),                                                                        //              (terminated)
		.uav_response             (),                                                                        //              (terminated)
		.av_response              (2'b00),                                                                   //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                    //              (terminated)
		.uav_writeresponsevalid   (),                                                                        //              (terminated)
		.av_writeresponserequest  (),                                                                        //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                     //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (22),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ch2_yn3_mu_s1_translator (
		.clk                      (clk_clk),                                                                  //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                       //                    reset.reset
		.uav_address              (ch2_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (ch2_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (ch2_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (ch2_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (ch2_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (ch2_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (ch2_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (ch2_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (ch2_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (ch2_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (ch2_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (ch2_yn3_mu_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (ch2_yn3_mu_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (ch2_yn3_mu_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (ch2_yn3_mu_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (ch2_yn3_mu_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                         //              (terminated)
		.av_begintransfer         (),                                                                         //              (terminated)
		.av_beginbursttransfer    (),                                                                         //              (terminated)
		.av_burstcount            (),                                                                         //              (terminated)
		.av_byteenable            (),                                                                         //              (terminated)
		.av_readdatavalid         (1'b0),                                                                     //              (terminated)
		.av_waitrequest           (1'b0),                                                                     //              (terminated)
		.av_writebyteenable       (),                                                                         //              (terminated)
		.av_lock                  (),                                                                         //              (terminated)
		.av_clken                 (),                                                                         //              (terminated)
		.uav_clken                (1'b0),                                                                     //              (terminated)
		.av_debugaccess           (),                                                                         //              (terminated)
		.av_outputenable          (),                                                                         //              (terminated)
		.uav_response             (),                                                                         //              (terminated)
		.av_response              (2'b00),                                                                    //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                     //              (terminated)
		.uav_writeresponsevalid   (),                                                                         //              (terminated)
		.av_writeresponserequest  (),                                                                         //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                      //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (22),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ch2_yn3_ml_s1_translator (
		.clk                      (clk_clk),                                                                  //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                       //                    reset.reset
		.uav_address              (ch2_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (ch2_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (ch2_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (ch2_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (ch2_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (ch2_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (ch2_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (ch2_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (ch2_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (ch2_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (ch2_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (ch2_yn3_ml_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (ch2_yn3_ml_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (ch2_yn3_ml_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (ch2_yn3_ml_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (ch2_yn3_ml_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                         //              (terminated)
		.av_begintransfer         (),                                                                         //              (terminated)
		.av_beginbursttransfer    (),                                                                         //              (terminated)
		.av_burstcount            (),                                                                         //              (terminated)
		.av_byteenable            (),                                                                         //              (terminated)
		.av_readdatavalid         (1'b0),                                                                     //              (terminated)
		.av_waitrequest           (1'b0),                                                                     //              (terminated)
		.av_writebyteenable       (),                                                                         //              (terminated)
		.av_lock                  (),                                                                         //              (terminated)
		.av_clken                 (),                                                                         //              (terminated)
		.uav_clken                (1'b0),                                                                     //              (terminated)
		.av_debugaccess           (),                                                                         //              (terminated)
		.av_outputenable          (),                                                                         //              (terminated)
		.uav_response             (),                                                                         //              (terminated)
		.av_response              (2'b00),                                                                    //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                     //              (terminated)
		.uav_writeresponsevalid   (),                                                                         //              (terminated)
		.av_writeresponserequest  (),                                                                         //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                      //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (22),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ch2_yn3_l_s1_translator (
		.clk                      (clk_clk),                                                                 //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                      //                    reset.reset
		.uav_address              (ch2_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (ch2_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (ch2_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (ch2_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (ch2_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (ch2_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (ch2_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (ch2_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (ch2_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (ch2_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (ch2_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (ch2_yn3_l_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (ch2_yn3_l_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (ch2_yn3_l_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (ch2_yn3_l_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (ch2_yn3_l_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                        //              (terminated)
		.av_begintransfer         (),                                                                        //              (terminated)
		.av_beginbursttransfer    (),                                                                        //              (terminated)
		.av_burstcount            (),                                                                        //              (terminated)
		.av_byteenable            (),                                                                        //              (terminated)
		.av_readdatavalid         (1'b0),                                                                    //              (terminated)
		.av_waitrequest           (1'b0),                                                                    //              (terminated)
		.av_writebyteenable       (),                                                                        //              (terminated)
		.av_lock                  (),                                                                        //              (terminated)
		.av_clken                 (),                                                                        //              (terminated)
		.uav_clken                (1'b0),                                                                    //              (terminated)
		.av_debugaccess           (),                                                                        //              (terminated)
		.av_outputenable          (),                                                                        //              (terminated)
		.uav_response             (),                                                                        //              (terminated)
		.av_response              (2'b00),                                                                   //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                    //              (terminated)
		.uav_writeresponsevalid   (),                                                                        //              (terminated)
		.av_writeresponserequest  (),                                                                        //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                     //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (22),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ch3_timer_rst_s1_translator (
		.clk                      (clk_clk),                                                                     //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                          //                    reset.reset
		.uav_address              (ch3_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (ch3_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (ch3_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (ch3_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (ch3_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (ch3_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (ch3_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (ch3_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (ch3_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (ch3_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (ch3_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (ch3_timer_rst_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (ch3_timer_rst_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (ch3_timer_rst_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (ch3_timer_rst_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (ch3_timer_rst_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                            //              (terminated)
		.av_begintransfer         (),                                                                            //              (terminated)
		.av_beginbursttransfer    (),                                                                            //              (terminated)
		.av_burstcount            (),                                                                            //              (terminated)
		.av_byteenable            (),                                                                            //              (terminated)
		.av_readdatavalid         (1'b0),                                                                        //              (terminated)
		.av_waitrequest           (1'b0),                                                                        //              (terminated)
		.av_writebyteenable       (),                                                                            //              (terminated)
		.av_lock                  (),                                                                            //              (terminated)
		.av_clken                 (),                                                                            //              (terminated)
		.uav_clken                (1'b0),                                                                        //              (terminated)
		.av_debugaccess           (),                                                                            //              (terminated)
		.av_outputenable          (),                                                                            //              (terminated)
		.uav_response             (),                                                                            //              (terminated)
		.av_response              (2'b00),                                                                       //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                        //              (terminated)
		.uav_writeresponsevalid   (),                                                                            //              (terminated)
		.av_writeresponserequest  (),                                                                            //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                         //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (22),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ch3_thresh_s1_translator (
		.clk                      (clk_clk),                                                                  //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                       //                    reset.reset
		.uav_address              (ch3_thresh_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (ch3_thresh_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (ch3_thresh_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (ch3_thresh_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (ch3_thresh_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (ch3_thresh_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (ch3_thresh_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (ch3_thresh_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (ch3_thresh_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (ch3_thresh_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (ch3_thresh_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (ch3_thresh_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (ch3_thresh_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (ch3_thresh_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (ch3_thresh_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (ch3_thresh_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                         //              (terminated)
		.av_begintransfer         (),                                                                         //              (terminated)
		.av_beginbursttransfer    (),                                                                         //              (terminated)
		.av_burstcount            (),                                                                         //              (terminated)
		.av_byteenable            (),                                                                         //              (terminated)
		.av_readdatavalid         (1'b0),                                                                     //              (terminated)
		.av_waitrequest           (1'b0),                                                                     //              (terminated)
		.av_writebyteenable       (),                                                                         //              (terminated)
		.av_lock                  (),                                                                         //              (terminated)
		.av_clken                 (),                                                                         //              (terminated)
		.uav_clken                (1'b0),                                                                     //              (terminated)
		.av_debugaccess           (),                                                                         //              (terminated)
		.av_outputenable          (),                                                                         //              (terminated)
		.uav_response             (),                                                                         //              (terminated)
		.av_response              (2'b00),                                                                    //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                     //              (terminated)
		.uav_writeresponsevalid   (),                                                                         //              (terminated)
		.av_writeresponserequest  (),                                                                         //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                      //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (22),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ch3_rd_peak_s1_translator (
		.clk                      (clk_clk),                                                                   //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                        //                    reset.reset
		.uav_address              (ch3_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (ch3_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (ch3_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (ch3_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (ch3_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (ch3_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (ch3_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (ch3_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (ch3_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (ch3_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (ch3_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (ch3_rd_peak_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (ch3_rd_peak_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (ch3_rd_peak_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (ch3_rd_peak_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (ch3_rd_peak_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                          //              (terminated)
		.av_begintransfer         (),                                                                          //              (terminated)
		.av_beginbursttransfer    (),                                                                          //              (terminated)
		.av_burstcount            (),                                                                          //              (terminated)
		.av_byteenable            (),                                                                          //              (terminated)
		.av_readdatavalid         (1'b0),                                                                      //              (terminated)
		.av_waitrequest           (1'b0),                                                                      //              (terminated)
		.av_writebyteenable       (),                                                                          //              (terminated)
		.av_lock                  (),                                                                          //              (terminated)
		.av_clken                 (),                                                                          //              (terminated)
		.uav_clken                (1'b0),                                                                      //              (terminated)
		.av_debugaccess           (),                                                                          //              (terminated)
		.av_outputenable          (),                                                                          //              (terminated)
		.uav_response             (),                                                                          //              (terminated)
		.av_response              (2'b00),                                                                     //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                      //              (terminated)
		.uav_writeresponsevalid   (),                                                                          //              (terminated)
		.av_writeresponserequest  (),                                                                          //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                       //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (22),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ch3_peak_found_s1_translator (
		.clk                      (clk_clk),                                                                      //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                           //                    reset.reset
		.uav_address              (ch3_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (ch3_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (ch3_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (ch3_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (ch3_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (ch3_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (ch3_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (ch3_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (ch3_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (ch3_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (ch3_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (ch3_peak_found_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (ch3_peak_found_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (ch3_peak_found_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (ch3_peak_found_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (ch3_peak_found_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                             //              (terminated)
		.av_begintransfer         (),                                                                             //              (terminated)
		.av_beginbursttransfer    (),                                                                             //              (terminated)
		.av_burstcount            (),                                                                             //              (terminated)
		.av_byteenable            (),                                                                             //              (terminated)
		.av_readdatavalid         (1'b0),                                                                         //              (terminated)
		.av_waitrequest           (1'b0),                                                                         //              (terminated)
		.av_writebyteenable       (),                                                                             //              (terminated)
		.av_lock                  (),                                                                             //              (terminated)
		.av_clken                 (),                                                                             //              (terminated)
		.uav_clken                (1'b0),                                                                         //              (terminated)
		.av_debugaccess           (),                                                                             //              (terminated)
		.av_outputenable          (),                                                                             //              (terminated)
		.uav_response             (),                                                                             //              (terminated)
		.av_response              (2'b00),                                                                        //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                         //              (terminated)
		.uav_writeresponsevalid   (),                                                                             //              (terminated)
		.av_writeresponserequest  (),                                                                             //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                          //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (22),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ch3_yn1_u_s1_translator (
		.clk                      (clk_clk),                                                                 //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                      //                    reset.reset
		.uav_address              (ch3_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (ch3_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (ch3_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (ch3_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (ch3_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (ch3_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (ch3_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (ch3_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (ch3_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (ch3_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (ch3_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (ch3_yn1_u_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (ch3_yn1_u_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (ch3_yn1_u_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (ch3_yn1_u_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (ch3_yn1_u_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                        //              (terminated)
		.av_begintransfer         (),                                                                        //              (terminated)
		.av_beginbursttransfer    (),                                                                        //              (terminated)
		.av_burstcount            (),                                                                        //              (terminated)
		.av_byteenable            (),                                                                        //              (terminated)
		.av_readdatavalid         (1'b0),                                                                    //              (terminated)
		.av_waitrequest           (1'b0),                                                                    //              (terminated)
		.av_writebyteenable       (),                                                                        //              (terminated)
		.av_lock                  (),                                                                        //              (terminated)
		.av_clken                 (),                                                                        //              (terminated)
		.uav_clken                (1'b0),                                                                    //              (terminated)
		.av_debugaccess           (),                                                                        //              (terminated)
		.av_outputenable          (),                                                                        //              (terminated)
		.uav_response             (),                                                                        //              (terminated)
		.av_response              (2'b00),                                                                   //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                    //              (terminated)
		.uav_writeresponsevalid   (),                                                                        //              (terminated)
		.av_writeresponserequest  (),                                                                        //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                     //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (22),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ch3_time_s1_translator (
		.clk                      (clk_clk),                                                                //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                     //                    reset.reset
		.uav_address              (ch3_time_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (ch3_time_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (ch3_time_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (ch3_time_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (ch3_time_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (ch3_time_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (ch3_time_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (ch3_time_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (ch3_time_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (ch3_time_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (ch3_time_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (ch3_time_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (ch3_time_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (ch3_time_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (ch3_time_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (ch3_time_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                       //              (terminated)
		.av_begintransfer         (),                                                                       //              (terminated)
		.av_beginbursttransfer    (),                                                                       //              (terminated)
		.av_burstcount            (),                                                                       //              (terminated)
		.av_byteenable            (),                                                                       //              (terminated)
		.av_readdatavalid         (1'b0),                                                                   //              (terminated)
		.av_waitrequest           (1'b0),                                                                   //              (terminated)
		.av_writebyteenable       (),                                                                       //              (terminated)
		.av_lock                  (),                                                                       //              (terminated)
		.av_clken                 (),                                                                       //              (terminated)
		.uav_clken                (1'b0),                                                                   //              (terminated)
		.av_debugaccess           (),                                                                       //              (terminated)
		.av_outputenable          (),                                                                       //              (terminated)
		.uav_response             (),                                                                       //              (terminated)
		.av_response              (2'b00),                                                                  //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                   //              (terminated)
		.uav_writeresponsevalid   (),                                                                       //              (terminated)
		.av_writeresponserequest  (),                                                                       //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                    //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (22),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ch3_yn3_l_s1_translator (
		.clk                      (clk_clk),                                                                 //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                      //                    reset.reset
		.uav_address              (ch3_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (ch3_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (ch3_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (ch3_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (ch3_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (ch3_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (ch3_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (ch3_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (ch3_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (ch3_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (ch3_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (ch3_yn3_l_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (ch3_yn3_l_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (ch3_yn3_l_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (ch3_yn3_l_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (ch3_yn3_l_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                        //              (terminated)
		.av_begintransfer         (),                                                                        //              (terminated)
		.av_beginbursttransfer    (),                                                                        //              (terminated)
		.av_burstcount            (),                                                                        //              (terminated)
		.av_byteenable            (),                                                                        //              (terminated)
		.av_readdatavalid         (1'b0),                                                                    //              (terminated)
		.av_waitrequest           (1'b0),                                                                    //              (terminated)
		.av_writebyteenable       (),                                                                        //              (terminated)
		.av_lock                  (),                                                                        //              (terminated)
		.av_clken                 (),                                                                        //              (terminated)
		.uav_clken                (1'b0),                                                                    //              (terminated)
		.av_debugaccess           (),                                                                        //              (terminated)
		.av_outputenable          (),                                                                        //              (terminated)
		.uav_response             (),                                                                        //              (terminated)
		.av_response              (2'b00),                                                                   //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                    //              (terminated)
		.uav_writeresponsevalid   (),                                                                        //              (terminated)
		.av_writeresponserequest  (),                                                                        //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                     //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (22),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ch3_yn3_ml_s1_translator (
		.clk                      (clk_clk),                                                                  //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                       //                    reset.reset
		.uav_address              (ch3_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (ch3_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (ch3_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (ch3_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (ch3_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (ch3_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (ch3_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (ch3_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (ch3_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (ch3_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (ch3_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (ch3_yn3_ml_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (ch3_yn3_ml_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (ch3_yn3_ml_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (ch3_yn3_ml_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (ch3_yn3_ml_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                         //              (terminated)
		.av_begintransfer         (),                                                                         //              (terminated)
		.av_beginbursttransfer    (),                                                                         //              (terminated)
		.av_burstcount            (),                                                                         //              (terminated)
		.av_byteenable            (),                                                                         //              (terminated)
		.av_readdatavalid         (1'b0),                                                                     //              (terminated)
		.av_waitrequest           (1'b0),                                                                     //              (terminated)
		.av_writebyteenable       (),                                                                         //              (terminated)
		.av_lock                  (),                                                                         //              (terminated)
		.av_clken                 (),                                                                         //              (terminated)
		.uav_clken                (1'b0),                                                                     //              (terminated)
		.av_debugaccess           (),                                                                         //              (terminated)
		.av_outputenable          (),                                                                         //              (terminated)
		.uav_response             (),                                                                         //              (terminated)
		.av_response              (2'b00),                                                                    //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                     //              (terminated)
		.uav_writeresponsevalid   (),                                                                         //              (terminated)
		.av_writeresponserequest  (),                                                                         //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                      //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (22),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ch3_yn3_mu_s1_translator (
		.clk                      (clk_clk),                                                                  //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                       //                    reset.reset
		.uav_address              (ch3_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (ch3_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (ch3_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (ch3_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (ch3_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (ch3_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (ch3_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (ch3_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (ch3_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (ch3_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (ch3_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (ch3_yn3_mu_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (ch3_yn3_mu_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (ch3_yn3_mu_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (ch3_yn3_mu_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (ch3_yn3_mu_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                         //              (terminated)
		.av_begintransfer         (),                                                                         //              (terminated)
		.av_beginbursttransfer    (),                                                                         //              (terminated)
		.av_burstcount            (),                                                                         //              (terminated)
		.av_byteenable            (),                                                                         //              (terminated)
		.av_readdatavalid         (1'b0),                                                                     //              (terminated)
		.av_waitrequest           (1'b0),                                                                     //              (terminated)
		.av_writebyteenable       (),                                                                         //              (terminated)
		.av_lock                  (),                                                                         //              (terminated)
		.av_clken                 (),                                                                         //              (terminated)
		.uav_clken                (1'b0),                                                                     //              (terminated)
		.av_debugaccess           (),                                                                         //              (terminated)
		.av_outputenable          (),                                                                         //              (terminated)
		.uav_response             (),                                                                         //              (terminated)
		.av_response              (2'b00),                                                                    //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                     //              (terminated)
		.uav_writeresponsevalid   (),                                                                         //              (terminated)
		.av_writeresponserequest  (),                                                                         //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                      //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (22),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ch3_yn3_u_s1_translator (
		.clk                      (clk_clk),                                                                 //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                      //                    reset.reset
		.uav_address              (ch3_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (ch3_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (ch3_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (ch3_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (ch3_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (ch3_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (ch3_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (ch3_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (ch3_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (ch3_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (ch3_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (ch3_yn3_u_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (ch3_yn3_u_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (ch3_yn3_u_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (ch3_yn3_u_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (ch3_yn3_u_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                        //              (terminated)
		.av_begintransfer         (),                                                                        //              (terminated)
		.av_beginbursttransfer    (),                                                                        //              (terminated)
		.av_burstcount            (),                                                                        //              (terminated)
		.av_byteenable            (),                                                                        //              (terminated)
		.av_readdatavalid         (1'b0),                                                                    //              (terminated)
		.av_waitrequest           (1'b0),                                                                    //              (terminated)
		.av_writebyteenable       (),                                                                        //              (terminated)
		.av_lock                  (),                                                                        //              (terminated)
		.av_clken                 (),                                                                        //              (terminated)
		.uav_clken                (1'b0),                                                                    //              (terminated)
		.av_debugaccess           (),                                                                        //              (terminated)
		.av_outputenable          (),                                                                        //              (terminated)
		.uav_response             (),                                                                        //              (terminated)
		.av_response              (2'b00),                                                                   //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                    //              (terminated)
		.uav_writeresponsevalid   (),                                                                        //              (terminated)
		.av_writeresponserequest  (),                                                                        //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                     //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (22),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ch3_yn2_l_s1_translator (
		.clk                      (clk_clk),                                                                 //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                      //                    reset.reset
		.uav_address              (ch3_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (ch3_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (ch3_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (ch3_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (ch3_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (ch3_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (ch3_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (ch3_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (ch3_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (ch3_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (ch3_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (ch3_yn2_l_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (ch3_yn2_l_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (ch3_yn2_l_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (ch3_yn2_l_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (ch3_yn2_l_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                        //              (terminated)
		.av_begintransfer         (),                                                                        //              (terminated)
		.av_beginbursttransfer    (),                                                                        //              (terminated)
		.av_burstcount            (),                                                                        //              (terminated)
		.av_byteenable            (),                                                                        //              (terminated)
		.av_readdatavalid         (1'b0),                                                                    //              (terminated)
		.av_waitrequest           (1'b0),                                                                    //              (terminated)
		.av_writebyteenable       (),                                                                        //              (terminated)
		.av_lock                  (),                                                                        //              (terminated)
		.av_clken                 (),                                                                        //              (terminated)
		.uav_clken                (1'b0),                                                                    //              (terminated)
		.av_debugaccess           (),                                                                        //              (terminated)
		.av_outputenable          (),                                                                        //              (terminated)
		.uav_response             (),                                                                        //              (terminated)
		.av_response              (2'b00),                                                                   //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                    //              (terminated)
		.uav_writeresponsevalid   (),                                                                        //              (terminated)
		.av_writeresponserequest  (),                                                                        //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                     //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (22),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ch3_yn2_ml_s1_translator (
		.clk                      (clk_clk),                                                                  //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                       //                    reset.reset
		.uav_address              (ch3_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (ch3_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (ch3_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (ch3_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (ch3_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (ch3_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (ch3_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (ch3_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (ch3_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (ch3_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (ch3_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (ch3_yn2_ml_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (ch3_yn2_ml_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (ch3_yn2_ml_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (ch3_yn2_ml_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (ch3_yn2_ml_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                         //              (terminated)
		.av_begintransfer         (),                                                                         //              (terminated)
		.av_beginbursttransfer    (),                                                                         //              (terminated)
		.av_burstcount            (),                                                                         //              (terminated)
		.av_byteenable            (),                                                                         //              (terminated)
		.av_readdatavalid         (1'b0),                                                                     //              (terminated)
		.av_waitrequest           (1'b0),                                                                     //              (terminated)
		.av_writebyteenable       (),                                                                         //              (terminated)
		.av_lock                  (),                                                                         //              (terminated)
		.av_clken                 (),                                                                         //              (terminated)
		.uav_clken                (1'b0),                                                                     //              (terminated)
		.av_debugaccess           (),                                                                         //              (terminated)
		.av_outputenable          (),                                                                         //              (terminated)
		.uav_response             (),                                                                         //              (terminated)
		.av_response              (2'b00),                                                                    //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                     //              (terminated)
		.uav_writeresponsevalid   (),                                                                         //              (terminated)
		.av_writeresponserequest  (),                                                                         //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                      //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (22),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ch3_yn2_mu_s1_translator (
		.clk                      (clk_clk),                                                                  //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                       //                    reset.reset
		.uav_address              (ch3_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (ch3_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (ch3_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (ch3_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (ch3_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (ch3_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (ch3_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (ch3_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (ch3_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (ch3_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (ch3_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (ch3_yn2_mu_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (ch3_yn2_mu_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (ch3_yn2_mu_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (ch3_yn2_mu_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (ch3_yn2_mu_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                         //              (terminated)
		.av_begintransfer         (),                                                                         //              (terminated)
		.av_beginbursttransfer    (),                                                                         //              (terminated)
		.av_burstcount            (),                                                                         //              (terminated)
		.av_byteenable            (),                                                                         //              (terminated)
		.av_readdatavalid         (1'b0),                                                                     //              (terminated)
		.av_waitrequest           (1'b0),                                                                     //              (terminated)
		.av_writebyteenable       (),                                                                         //              (terminated)
		.av_lock                  (),                                                                         //              (terminated)
		.av_clken                 (),                                                                         //              (terminated)
		.uav_clken                (1'b0),                                                                     //              (terminated)
		.av_debugaccess           (),                                                                         //              (terminated)
		.av_outputenable          (),                                                                         //              (terminated)
		.uav_response             (),                                                                         //              (terminated)
		.av_response              (2'b00),                                                                    //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                     //              (terminated)
		.uav_writeresponsevalid   (),                                                                         //              (terminated)
		.av_writeresponserequest  (),                                                                         //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                      //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (22),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ch3_yn2_u_s1_translator (
		.clk                      (clk_clk),                                                                 //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                      //                    reset.reset
		.uav_address              (ch3_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (ch3_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (ch3_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (ch3_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (ch3_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (ch3_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (ch3_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (ch3_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (ch3_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (ch3_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (ch3_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (ch3_yn2_u_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (ch3_yn2_u_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (ch3_yn2_u_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (ch3_yn2_u_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (ch3_yn2_u_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                        //              (terminated)
		.av_begintransfer         (),                                                                        //              (terminated)
		.av_beginbursttransfer    (),                                                                        //              (terminated)
		.av_burstcount            (),                                                                        //              (terminated)
		.av_byteenable            (),                                                                        //              (terminated)
		.av_readdatavalid         (1'b0),                                                                    //              (terminated)
		.av_waitrequest           (1'b0),                                                                    //              (terminated)
		.av_writebyteenable       (),                                                                        //              (terminated)
		.av_lock                  (),                                                                        //              (terminated)
		.av_clken                 (),                                                                        //              (terminated)
		.uav_clken                (1'b0),                                                                    //              (terminated)
		.av_debugaccess           (),                                                                        //              (terminated)
		.av_outputenable          (),                                                                        //              (terminated)
		.uav_response             (),                                                                        //              (terminated)
		.av_response              (2'b00),                                                                   //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                    //              (terminated)
		.uav_writeresponsevalid   (),                                                                        //              (terminated)
		.av_writeresponserequest  (),                                                                        //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                     //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (22),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ch3_yn1_l_s1_translator (
		.clk                      (clk_clk),                                                                 //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                      //                    reset.reset
		.uav_address              (ch3_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (ch3_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (ch3_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (ch3_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (ch3_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (ch3_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (ch3_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (ch3_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (ch3_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (ch3_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (ch3_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (ch3_yn1_l_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (ch3_yn1_l_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (ch3_yn1_l_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (ch3_yn1_l_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (ch3_yn1_l_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                        //              (terminated)
		.av_begintransfer         (),                                                                        //              (terminated)
		.av_beginbursttransfer    (),                                                                        //              (terminated)
		.av_burstcount            (),                                                                        //              (terminated)
		.av_byteenable            (),                                                                        //              (terminated)
		.av_readdatavalid         (1'b0),                                                                    //              (terminated)
		.av_waitrequest           (1'b0),                                                                    //              (terminated)
		.av_writebyteenable       (),                                                                        //              (terminated)
		.av_lock                  (),                                                                        //              (terminated)
		.av_clken                 (),                                                                        //              (terminated)
		.uav_clken                (1'b0),                                                                    //              (terminated)
		.av_debugaccess           (),                                                                        //              (terminated)
		.av_outputenable          (),                                                                        //              (terminated)
		.uav_response             (),                                                                        //              (terminated)
		.av_response              (2'b00),                                                                   //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                    //              (terminated)
		.uav_writeresponsevalid   (),                                                                        //              (terminated)
		.av_writeresponserequest  (),                                                                        //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                     //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (22),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ch3_yn1_mu_s1_translator (
		.clk                      (clk_clk),                                                                  //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                       //                    reset.reset
		.uav_address              (ch3_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (ch3_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (ch3_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (ch3_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (ch3_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (ch3_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (ch3_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (ch3_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (ch3_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (ch3_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (ch3_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (ch3_yn1_mu_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (ch3_yn1_mu_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (ch3_yn1_mu_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (ch3_yn1_mu_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (ch3_yn1_mu_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                         //              (terminated)
		.av_begintransfer         (),                                                                         //              (terminated)
		.av_beginbursttransfer    (),                                                                         //              (terminated)
		.av_burstcount            (),                                                                         //              (terminated)
		.av_byteenable            (),                                                                         //              (terminated)
		.av_readdatavalid         (1'b0),                                                                     //              (terminated)
		.av_waitrequest           (1'b0),                                                                     //              (terminated)
		.av_writebyteenable       (),                                                                         //              (terminated)
		.av_lock                  (),                                                                         //              (terminated)
		.av_clken                 (),                                                                         //              (terminated)
		.uav_clken                (1'b0),                                                                     //              (terminated)
		.av_debugaccess           (),                                                                         //              (terminated)
		.av_outputenable          (),                                                                         //              (terminated)
		.uav_response             (),                                                                         //              (terminated)
		.av_response              (2'b00),                                                                    //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                     //              (terminated)
		.uav_writeresponsevalid   (),                                                                         //              (terminated)
		.av_writeresponserequest  (),                                                                         //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                      //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (22),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ch3_yn1_ml_s1_translator (
		.clk                      (clk_clk),                                                                  //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                       //                    reset.reset
		.uav_address              (ch3_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (ch3_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (ch3_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (ch3_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (ch3_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (ch3_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (ch3_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (ch3_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (ch3_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (ch3_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (ch3_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (ch3_yn1_ml_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (ch3_yn1_ml_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (ch3_yn1_ml_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (ch3_yn1_ml_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (ch3_yn1_ml_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                         //              (terminated)
		.av_begintransfer         (),                                                                         //              (terminated)
		.av_beginbursttransfer    (),                                                                         //              (terminated)
		.av_burstcount            (),                                                                         //              (terminated)
		.av_byteenable            (),                                                                         //              (terminated)
		.av_readdatavalid         (1'b0),                                                                     //              (terminated)
		.av_waitrequest           (1'b0),                                                                     //              (terminated)
		.av_writebyteenable       (),                                                                         //              (terminated)
		.av_lock                  (),                                                                         //              (terminated)
		.av_clken                 (),                                                                         //              (terminated)
		.uav_clken                (1'b0),                                                                     //              (terminated)
		.av_debugaccess           (),                                                                         //              (terminated)
		.av_outputenable          (),                                                                         //              (terminated)
		.uav_response             (),                                                                         //              (terminated)
		.av_response              (2'b00),                                                                    //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                     //              (terminated)
		.uav_writeresponsevalid   (),                                                                         //              (terminated)
		.av_writeresponserequest  (),                                                                         //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                      //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (22),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ch4_timer_rst_s1_translator (
		.clk                      (clk_clk),                                                                     //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                          //                    reset.reset
		.uav_address              (ch4_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (ch4_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (ch4_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (ch4_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (ch4_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (ch4_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (ch4_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (ch4_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (ch4_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (ch4_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (ch4_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (ch4_timer_rst_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (ch4_timer_rst_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (ch4_timer_rst_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (ch4_timer_rst_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (ch4_timer_rst_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                            //              (terminated)
		.av_begintransfer         (),                                                                            //              (terminated)
		.av_beginbursttransfer    (),                                                                            //              (terminated)
		.av_burstcount            (),                                                                            //              (terminated)
		.av_byteenable            (),                                                                            //              (terminated)
		.av_readdatavalid         (1'b0),                                                                        //              (terminated)
		.av_waitrequest           (1'b0),                                                                        //              (terminated)
		.av_writebyteenable       (),                                                                            //              (terminated)
		.av_lock                  (),                                                                            //              (terminated)
		.av_clken                 (),                                                                            //              (terminated)
		.uav_clken                (1'b0),                                                                        //              (terminated)
		.av_debugaccess           (),                                                                            //              (terminated)
		.av_outputenable          (),                                                                            //              (terminated)
		.uav_response             (),                                                                            //              (terminated)
		.av_response              (2'b00),                                                                       //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                        //              (terminated)
		.uav_writeresponsevalid   (),                                                                            //              (terminated)
		.av_writeresponserequest  (),                                                                            //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                         //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (22),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ch4_thresh_s1_translator (
		.clk                      (clk_clk),                                                                  //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                       //                    reset.reset
		.uav_address              (ch4_thresh_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (ch4_thresh_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (ch4_thresh_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (ch4_thresh_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (ch4_thresh_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (ch4_thresh_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (ch4_thresh_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (ch4_thresh_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (ch4_thresh_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (ch4_thresh_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (ch4_thresh_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (ch4_thresh_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (ch4_thresh_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (ch4_thresh_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (ch4_thresh_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (ch4_thresh_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                         //              (terminated)
		.av_begintransfer         (),                                                                         //              (terminated)
		.av_beginbursttransfer    (),                                                                         //              (terminated)
		.av_burstcount            (),                                                                         //              (terminated)
		.av_byteenable            (),                                                                         //              (terminated)
		.av_readdatavalid         (1'b0),                                                                     //              (terminated)
		.av_waitrequest           (1'b0),                                                                     //              (terminated)
		.av_writebyteenable       (),                                                                         //              (terminated)
		.av_lock                  (),                                                                         //              (terminated)
		.av_clken                 (),                                                                         //              (terminated)
		.uav_clken                (1'b0),                                                                     //              (terminated)
		.av_debugaccess           (),                                                                         //              (terminated)
		.av_outputenable          (),                                                                         //              (terminated)
		.uav_response             (),                                                                         //              (terminated)
		.av_response              (2'b00),                                                                    //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                     //              (terminated)
		.uav_writeresponsevalid   (),                                                                         //              (terminated)
		.av_writeresponserequest  (),                                                                         //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                      //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (22),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ch4_rd_peak_s1_translator (
		.clk                      (clk_clk),                                                                   //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                        //                    reset.reset
		.uav_address              (ch4_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (ch4_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (ch4_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (ch4_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (ch4_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (ch4_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (ch4_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (ch4_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (ch4_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (ch4_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (ch4_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (ch4_rd_peak_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (ch4_rd_peak_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (ch4_rd_peak_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (ch4_rd_peak_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (ch4_rd_peak_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                          //              (terminated)
		.av_begintransfer         (),                                                                          //              (terminated)
		.av_beginbursttransfer    (),                                                                          //              (terminated)
		.av_burstcount            (),                                                                          //              (terminated)
		.av_byteenable            (),                                                                          //              (terminated)
		.av_readdatavalid         (1'b0),                                                                      //              (terminated)
		.av_waitrequest           (1'b0),                                                                      //              (terminated)
		.av_writebyteenable       (),                                                                          //              (terminated)
		.av_lock                  (),                                                                          //              (terminated)
		.av_clken                 (),                                                                          //              (terminated)
		.uav_clken                (1'b0),                                                                      //              (terminated)
		.av_debugaccess           (),                                                                          //              (terminated)
		.av_outputenable          (),                                                                          //              (terminated)
		.uav_response             (),                                                                          //              (terminated)
		.av_response              (2'b00),                                                                     //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                      //              (terminated)
		.uav_writeresponsevalid   (),                                                                          //              (terminated)
		.av_writeresponserequest  (),                                                                          //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                       //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (22),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ch4_peak_found_s1_translator (
		.clk                      (clk_clk),                                                                      //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                           //                    reset.reset
		.uav_address              (ch4_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (ch4_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (ch4_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (ch4_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (ch4_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (ch4_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (ch4_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (ch4_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (ch4_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (ch4_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (ch4_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (ch4_peak_found_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (ch4_peak_found_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (ch4_peak_found_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (ch4_peak_found_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (ch4_peak_found_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                             //              (terminated)
		.av_begintransfer         (),                                                                             //              (terminated)
		.av_beginbursttransfer    (),                                                                             //              (terminated)
		.av_burstcount            (),                                                                             //              (terminated)
		.av_byteenable            (),                                                                             //              (terminated)
		.av_readdatavalid         (1'b0),                                                                         //              (terminated)
		.av_waitrequest           (1'b0),                                                                         //              (terminated)
		.av_writebyteenable       (),                                                                             //              (terminated)
		.av_lock                  (),                                                                             //              (terminated)
		.av_clken                 (),                                                                             //              (terminated)
		.uav_clken                (1'b0),                                                                         //              (terminated)
		.av_debugaccess           (),                                                                             //              (terminated)
		.av_outputenable          (),                                                                             //              (terminated)
		.uav_response             (),                                                                             //              (terminated)
		.av_response              (2'b00),                                                                        //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                         //              (terminated)
		.uav_writeresponsevalid   (),                                                                             //              (terminated)
		.av_writeresponserequest  (),                                                                             //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                          //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (22),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ch4_time_s1_translator (
		.clk                      (clk_clk),                                                                //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                     //                    reset.reset
		.uav_address              (ch4_time_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (ch4_time_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (ch4_time_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (ch4_time_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (ch4_time_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (ch4_time_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (ch4_time_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (ch4_time_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (ch4_time_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (ch4_time_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (ch4_time_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (ch4_time_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (ch4_time_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (ch4_time_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (ch4_time_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (ch4_time_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                       //              (terminated)
		.av_begintransfer         (),                                                                       //              (terminated)
		.av_beginbursttransfer    (),                                                                       //              (terminated)
		.av_burstcount            (),                                                                       //              (terminated)
		.av_byteenable            (),                                                                       //              (terminated)
		.av_readdatavalid         (1'b0),                                                                   //              (terminated)
		.av_waitrequest           (1'b0),                                                                   //              (terminated)
		.av_writebyteenable       (),                                                                       //              (terminated)
		.av_lock                  (),                                                                       //              (terminated)
		.av_clken                 (),                                                                       //              (terminated)
		.uav_clken                (1'b0),                                                                   //              (terminated)
		.av_debugaccess           (),                                                                       //              (terminated)
		.av_outputenable          (),                                                                       //              (terminated)
		.uav_response             (),                                                                       //              (terminated)
		.av_response              (2'b00),                                                                  //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                   //              (terminated)
		.uav_writeresponsevalid   (),                                                                       //              (terminated)
		.av_writeresponserequest  (),                                                                       //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                    //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (22),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ch4_yn1_u_s1_translator (
		.clk                      (clk_clk),                                                                 //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                      //                    reset.reset
		.uav_address              (ch4_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (ch4_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (ch4_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (ch4_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (ch4_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (ch4_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (ch4_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (ch4_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (ch4_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (ch4_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (ch4_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (ch4_yn1_u_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (ch4_yn1_u_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (ch4_yn1_u_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (ch4_yn1_u_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (ch4_yn1_u_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                        //              (terminated)
		.av_begintransfer         (),                                                                        //              (terminated)
		.av_beginbursttransfer    (),                                                                        //              (terminated)
		.av_burstcount            (),                                                                        //              (terminated)
		.av_byteenable            (),                                                                        //              (terminated)
		.av_readdatavalid         (1'b0),                                                                    //              (terminated)
		.av_waitrequest           (1'b0),                                                                    //              (terminated)
		.av_writebyteenable       (),                                                                        //              (terminated)
		.av_lock                  (),                                                                        //              (terminated)
		.av_clken                 (),                                                                        //              (terminated)
		.uav_clken                (1'b0),                                                                    //              (terminated)
		.av_debugaccess           (),                                                                        //              (terminated)
		.av_outputenable          (),                                                                        //              (terminated)
		.uav_response             (),                                                                        //              (terminated)
		.av_response              (2'b00),                                                                   //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                    //              (terminated)
		.uav_writeresponsevalid   (),                                                                        //              (terminated)
		.av_writeresponserequest  (),                                                                        //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                     //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (22),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ch4_yn1_mu_s1_translator (
		.clk                      (clk_clk),                                                                  //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                       //                    reset.reset
		.uav_address              (ch4_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (ch4_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (ch4_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (ch4_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (ch4_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (ch4_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (ch4_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (ch4_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (ch4_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (ch4_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (ch4_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (ch4_yn1_mu_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (ch4_yn1_mu_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (ch4_yn1_mu_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (ch4_yn1_mu_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (ch4_yn1_mu_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                         //              (terminated)
		.av_begintransfer         (),                                                                         //              (terminated)
		.av_beginbursttransfer    (),                                                                         //              (terminated)
		.av_burstcount            (),                                                                         //              (terminated)
		.av_byteenable            (),                                                                         //              (terminated)
		.av_readdatavalid         (1'b0),                                                                     //              (terminated)
		.av_waitrequest           (1'b0),                                                                     //              (terminated)
		.av_writebyteenable       (),                                                                         //              (terminated)
		.av_lock                  (),                                                                         //              (terminated)
		.av_clken                 (),                                                                         //              (terminated)
		.uav_clken                (1'b0),                                                                     //              (terminated)
		.av_debugaccess           (),                                                                         //              (terminated)
		.av_outputenable          (),                                                                         //              (terminated)
		.uav_response             (),                                                                         //              (terminated)
		.av_response              (2'b00),                                                                    //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                     //              (terminated)
		.uav_writeresponsevalid   (),                                                                         //              (terminated)
		.av_writeresponserequest  (),                                                                         //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                      //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (22),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ch4_yn1_ml_s1_translator (
		.clk                      (clk_clk),                                                                  //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                       //                    reset.reset
		.uav_address              (ch4_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (ch4_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (ch4_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (ch4_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (ch4_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (ch4_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (ch4_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (ch4_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (ch4_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (ch4_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (ch4_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (ch4_yn1_ml_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (ch4_yn1_ml_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (ch4_yn1_ml_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (ch4_yn1_ml_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (ch4_yn1_ml_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                         //              (terminated)
		.av_begintransfer         (),                                                                         //              (terminated)
		.av_beginbursttransfer    (),                                                                         //              (terminated)
		.av_burstcount            (),                                                                         //              (terminated)
		.av_byteenable            (),                                                                         //              (terminated)
		.av_readdatavalid         (1'b0),                                                                     //              (terminated)
		.av_waitrequest           (1'b0),                                                                     //              (terminated)
		.av_writebyteenable       (),                                                                         //              (terminated)
		.av_lock                  (),                                                                         //              (terminated)
		.av_clken                 (),                                                                         //              (terminated)
		.uav_clken                (1'b0),                                                                     //              (terminated)
		.av_debugaccess           (),                                                                         //              (terminated)
		.av_outputenable          (),                                                                         //              (terminated)
		.uav_response             (),                                                                         //              (terminated)
		.av_response              (2'b00),                                                                    //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                     //              (terminated)
		.uav_writeresponsevalid   (),                                                                         //              (terminated)
		.av_writeresponserequest  (),                                                                         //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                      //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (22),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ch4_yn1_l_s1_translator (
		.clk                      (clk_clk),                                                                 //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                      //                    reset.reset
		.uav_address              (ch4_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (ch4_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (ch4_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (ch4_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (ch4_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (ch4_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (ch4_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (ch4_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (ch4_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (ch4_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (ch4_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (ch4_yn1_l_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (ch4_yn1_l_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (ch4_yn1_l_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (ch4_yn1_l_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (ch4_yn1_l_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                        //              (terminated)
		.av_begintransfer         (),                                                                        //              (terminated)
		.av_beginbursttransfer    (),                                                                        //              (terminated)
		.av_burstcount            (),                                                                        //              (terminated)
		.av_byteenable            (),                                                                        //              (terminated)
		.av_readdatavalid         (1'b0),                                                                    //              (terminated)
		.av_waitrequest           (1'b0),                                                                    //              (terminated)
		.av_writebyteenable       (),                                                                        //              (terminated)
		.av_lock                  (),                                                                        //              (terminated)
		.av_clken                 (),                                                                        //              (terminated)
		.uav_clken                (1'b0),                                                                    //              (terminated)
		.av_debugaccess           (),                                                                        //              (terminated)
		.av_outputenable          (),                                                                        //              (terminated)
		.uav_response             (),                                                                        //              (terminated)
		.av_response              (2'b00),                                                                   //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                    //              (terminated)
		.uav_writeresponsevalid   (),                                                                        //              (terminated)
		.av_writeresponserequest  (),                                                                        //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                     //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (22),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ch4_yn2_u_s1_translator (
		.clk                      (clk_clk),                                                                 //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                      //                    reset.reset
		.uav_address              (ch4_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (ch4_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (ch4_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (ch4_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (ch4_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (ch4_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (ch4_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (ch4_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (ch4_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (ch4_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (ch4_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (ch4_yn2_u_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (ch4_yn2_u_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (ch4_yn2_u_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (ch4_yn2_u_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (ch4_yn2_u_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                        //              (terminated)
		.av_begintransfer         (),                                                                        //              (terminated)
		.av_beginbursttransfer    (),                                                                        //              (terminated)
		.av_burstcount            (),                                                                        //              (terminated)
		.av_byteenable            (),                                                                        //              (terminated)
		.av_readdatavalid         (1'b0),                                                                    //              (terminated)
		.av_waitrequest           (1'b0),                                                                    //              (terminated)
		.av_writebyteenable       (),                                                                        //              (terminated)
		.av_lock                  (),                                                                        //              (terminated)
		.av_clken                 (),                                                                        //              (terminated)
		.uav_clken                (1'b0),                                                                    //              (terminated)
		.av_debugaccess           (),                                                                        //              (terminated)
		.av_outputenable          (),                                                                        //              (terminated)
		.uav_response             (),                                                                        //              (terminated)
		.av_response              (2'b00),                                                                   //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                    //              (terminated)
		.uav_writeresponsevalid   (),                                                                        //              (terminated)
		.av_writeresponserequest  (),                                                                        //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                     //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (22),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ch4_yn2_mu_s1_translator (
		.clk                      (clk_clk),                                                                  //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                       //                    reset.reset
		.uav_address              (ch4_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (ch4_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (ch4_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (ch4_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (ch4_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (ch4_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (ch4_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (ch4_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (ch4_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (ch4_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (ch4_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (ch4_yn2_mu_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (ch4_yn2_mu_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (ch4_yn2_mu_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (ch4_yn2_mu_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (ch4_yn2_mu_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                         //              (terminated)
		.av_begintransfer         (),                                                                         //              (terminated)
		.av_beginbursttransfer    (),                                                                         //              (terminated)
		.av_burstcount            (),                                                                         //              (terminated)
		.av_byteenable            (),                                                                         //              (terminated)
		.av_readdatavalid         (1'b0),                                                                     //              (terminated)
		.av_waitrequest           (1'b0),                                                                     //              (terminated)
		.av_writebyteenable       (),                                                                         //              (terminated)
		.av_lock                  (),                                                                         //              (terminated)
		.av_clken                 (),                                                                         //              (terminated)
		.uav_clken                (1'b0),                                                                     //              (terminated)
		.av_debugaccess           (),                                                                         //              (terminated)
		.av_outputenable          (),                                                                         //              (terminated)
		.uav_response             (),                                                                         //              (terminated)
		.av_response              (2'b00),                                                                    //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                     //              (terminated)
		.uav_writeresponsevalid   (),                                                                         //              (terminated)
		.av_writeresponserequest  (),                                                                         //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                      //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (22),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ch4_yn2_ml_s1_translator (
		.clk                      (clk_clk),                                                                  //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                       //                    reset.reset
		.uav_address              (ch4_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (ch4_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (ch4_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (ch4_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (ch4_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (ch4_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (ch4_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (ch4_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (ch4_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (ch4_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (ch4_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (ch4_yn2_ml_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (ch4_yn2_ml_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (ch4_yn2_ml_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (ch4_yn2_ml_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (ch4_yn2_ml_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                         //              (terminated)
		.av_begintransfer         (),                                                                         //              (terminated)
		.av_beginbursttransfer    (),                                                                         //              (terminated)
		.av_burstcount            (),                                                                         //              (terminated)
		.av_byteenable            (),                                                                         //              (terminated)
		.av_readdatavalid         (1'b0),                                                                     //              (terminated)
		.av_waitrequest           (1'b0),                                                                     //              (terminated)
		.av_writebyteenable       (),                                                                         //              (terminated)
		.av_lock                  (),                                                                         //              (terminated)
		.av_clken                 (),                                                                         //              (terminated)
		.uav_clken                (1'b0),                                                                     //              (terminated)
		.av_debugaccess           (),                                                                         //              (terminated)
		.av_outputenable          (),                                                                         //              (terminated)
		.uav_response             (),                                                                         //              (terminated)
		.av_response              (2'b00),                                                                    //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                     //              (terminated)
		.uav_writeresponsevalid   (),                                                                         //              (terminated)
		.av_writeresponserequest  (),                                                                         //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                      //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (22),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ch4_yn2_l_s1_translator (
		.clk                      (clk_clk),                                                                 //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                      //                    reset.reset
		.uav_address              (ch4_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (ch4_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (ch4_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (ch4_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (ch4_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (ch4_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (ch4_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (ch4_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (ch4_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (ch4_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (ch4_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (ch4_yn2_l_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (ch4_yn2_l_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (ch4_yn2_l_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (ch4_yn2_l_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (ch4_yn2_l_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                        //              (terminated)
		.av_begintransfer         (),                                                                        //              (terminated)
		.av_beginbursttransfer    (),                                                                        //              (terminated)
		.av_burstcount            (),                                                                        //              (terminated)
		.av_byteenable            (),                                                                        //              (terminated)
		.av_readdatavalid         (1'b0),                                                                    //              (terminated)
		.av_waitrequest           (1'b0),                                                                    //              (terminated)
		.av_writebyteenable       (),                                                                        //              (terminated)
		.av_lock                  (),                                                                        //              (terminated)
		.av_clken                 (),                                                                        //              (terminated)
		.uav_clken                (1'b0),                                                                    //              (terminated)
		.av_debugaccess           (),                                                                        //              (terminated)
		.av_outputenable          (),                                                                        //              (terminated)
		.uav_response             (),                                                                        //              (terminated)
		.av_response              (2'b00),                                                                   //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                    //              (terminated)
		.uav_writeresponsevalid   (),                                                                        //              (terminated)
		.av_writeresponserequest  (),                                                                        //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                     //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (22),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ch4_yn3_u_s1_translator (
		.clk                      (clk_clk),                                                                 //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                      //                    reset.reset
		.uav_address              (ch4_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (ch4_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (ch4_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (ch4_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (ch4_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (ch4_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (ch4_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (ch4_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (ch4_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (ch4_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (ch4_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (ch4_yn3_u_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (ch4_yn3_u_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (ch4_yn3_u_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (ch4_yn3_u_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (ch4_yn3_u_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                        //              (terminated)
		.av_begintransfer         (),                                                                        //              (terminated)
		.av_beginbursttransfer    (),                                                                        //              (terminated)
		.av_burstcount            (),                                                                        //              (terminated)
		.av_byteenable            (),                                                                        //              (terminated)
		.av_readdatavalid         (1'b0),                                                                    //              (terminated)
		.av_waitrequest           (1'b0),                                                                    //              (terminated)
		.av_writebyteenable       (),                                                                        //              (terminated)
		.av_lock                  (),                                                                        //              (terminated)
		.av_clken                 (),                                                                        //              (terminated)
		.uav_clken                (1'b0),                                                                    //              (terminated)
		.av_debugaccess           (),                                                                        //              (terminated)
		.av_outputenable          (),                                                                        //              (terminated)
		.uav_response             (),                                                                        //              (terminated)
		.av_response              (2'b00),                                                                   //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                    //              (terminated)
		.uav_writeresponsevalid   (),                                                                        //              (terminated)
		.av_writeresponserequest  (),                                                                        //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                     //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (22),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ch4_yn3_mu_s1_translator (
		.clk                      (clk_clk),                                                                  //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                       //                    reset.reset
		.uav_address              (ch4_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (ch4_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (ch4_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (ch4_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (ch4_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (ch4_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (ch4_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (ch4_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (ch4_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (ch4_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (ch4_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (ch4_yn3_mu_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (ch4_yn3_mu_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (ch4_yn3_mu_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (ch4_yn3_mu_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (ch4_yn3_mu_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                         //              (terminated)
		.av_begintransfer         (),                                                                         //              (terminated)
		.av_beginbursttransfer    (),                                                                         //              (terminated)
		.av_burstcount            (),                                                                         //              (terminated)
		.av_byteenable            (),                                                                         //              (terminated)
		.av_readdatavalid         (1'b0),                                                                     //              (terminated)
		.av_waitrequest           (1'b0),                                                                     //              (terminated)
		.av_writebyteenable       (),                                                                         //              (terminated)
		.av_lock                  (),                                                                         //              (terminated)
		.av_clken                 (),                                                                         //              (terminated)
		.uav_clken                (1'b0),                                                                     //              (terminated)
		.av_debugaccess           (),                                                                         //              (terminated)
		.av_outputenable          (),                                                                         //              (terminated)
		.uav_response             (),                                                                         //              (terminated)
		.av_response              (2'b00),                                                                    //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                     //              (terminated)
		.uav_writeresponsevalid   (),                                                                         //              (terminated)
		.av_writeresponserequest  (),                                                                         //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                      //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (22),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ch4_yn3_ml_s1_translator (
		.clk                      (clk_clk),                                                                  //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                       //                    reset.reset
		.uav_address              (ch4_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (ch4_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (ch4_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (ch4_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (ch4_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (ch4_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (ch4_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (ch4_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (ch4_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (ch4_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (ch4_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (ch4_yn3_ml_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (ch4_yn3_ml_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (ch4_yn3_ml_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (ch4_yn3_ml_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (ch4_yn3_ml_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                         //              (terminated)
		.av_begintransfer         (),                                                                         //              (terminated)
		.av_beginbursttransfer    (),                                                                         //              (terminated)
		.av_burstcount            (),                                                                         //              (terminated)
		.av_byteenable            (),                                                                         //              (terminated)
		.av_readdatavalid         (1'b0),                                                                     //              (terminated)
		.av_waitrequest           (1'b0),                                                                     //              (terminated)
		.av_writebyteenable       (),                                                                         //              (terminated)
		.av_lock                  (),                                                                         //              (terminated)
		.av_clken                 (),                                                                         //              (terminated)
		.uav_clken                (1'b0),                                                                     //              (terminated)
		.av_debugaccess           (),                                                                         //              (terminated)
		.av_outputenable          (),                                                                         //              (terminated)
		.uav_response             (),                                                                         //              (terminated)
		.av_response              (2'b00),                                                                    //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                     //              (terminated)
		.uav_writeresponsevalid   (),                                                                         //              (terminated)
		.av_writeresponserequest  (),                                                                         //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                      //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (22),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ch4_yn3_l_s1_translator (
		.clk                      (clk_clk),                                                                 //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                      //                    reset.reset
		.uav_address              (ch4_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (ch4_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (ch4_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (ch4_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (ch4_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (ch4_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (ch4_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (ch4_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (ch4_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (ch4_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (ch4_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (ch4_yn3_l_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (ch4_yn3_l_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (ch4_yn3_l_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (ch4_yn3_l_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (ch4_yn3_l_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                        //              (terminated)
		.av_begintransfer         (),                                                                        //              (terminated)
		.av_beginbursttransfer    (),                                                                        //              (terminated)
		.av_burstcount            (),                                                                        //              (terminated)
		.av_byteenable            (),                                                                        //              (terminated)
		.av_readdatavalid         (1'b0),                                                                    //              (terminated)
		.av_waitrequest           (1'b0),                                                                    //              (terminated)
		.av_writebyteenable       (),                                                                        //              (terminated)
		.av_lock                  (),                                                                        //              (terminated)
		.av_clken                 (),                                                                        //              (terminated)
		.uav_clken                (1'b0),                                                                    //              (terminated)
		.av_debugaccess           (),                                                                        //              (terminated)
		.av_outputenable          (),                                                                        //              (terminated)
		.uav_response             (),                                                                        //              (terminated)
		.av_response              (2'b00),                                                                   //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                    //              (terminated)
		.uav_writeresponsevalid   (),                                                                        //              (terminated)
		.av_writeresponserequest  (),                                                                        //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                     //              (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_BEGIN_BURST           (77),
		.PKT_BURSTWRAP_H           (69),
		.PKT_BURSTWRAP_L           (67),
		.PKT_BURST_SIZE_H          (72),
		.PKT_BURST_SIZE_L          (70),
		.PKT_BURST_TYPE_H          (74),
		.PKT_BURST_TYPE_L          (73),
		.PKT_BYTE_CNT_H            (66),
		.PKT_BYTE_CNT_L            (64),
		.PKT_ADDR_H                (57),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (58),
		.PKT_TRANS_POSTED          (59),
		.PKT_TRANS_WRITE           (60),
		.PKT_TRANS_READ            (61),
		.PKT_TRANS_LOCK            (62),
		.PKT_TRANS_EXCLUSIVE       (63),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (85),
		.PKT_SRC_ID_L              (79),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (86),
		.PKT_THREAD_ID_H           (93),
		.PKT_THREAD_ID_L           (93),
		.PKT_CACHE_H               (100),
		.PKT_CACHE_L               (97),
		.PKT_DATA_SIDEBAND_H       (76),
		.PKT_DATA_SIDEBAND_L       (76),
		.PKT_QOS_H                 (78),
		.PKT_QOS_L                 (78),
		.PKT_ADDR_SIDEBAND_H       (75),
		.PKT_ADDR_SIDEBAND_L       (75),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.ST_DATA_W                 (103),
		.ST_CHANNEL_W              (99),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (1),
		.BURSTWRAP_VALUE           (3),
		.CACHE_VALUE               (0),
		.SECURE_ACCESS_BIT         (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) nios_cpu_instruction_master_translator_avalon_universal_master_0_agent (
		.clk                     (clk_clk),                                                                                 //       clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                          // clk_reset.reset
		.av_address              (nios_cpu_instruction_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write                (nios_cpu_instruction_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read                 (nios_cpu_instruction_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata            (nios_cpu_instruction_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata             (nios_cpu_instruction_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest          (nios_cpu_instruction_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid        (nios_cpu_instruction_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable           (nios_cpu_instruction_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount           (nios_cpu_instruction_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess          (nios_cpu_instruction_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock                 (nios_cpu_instruction_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid                (nios_cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data                 (nios_cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket        (nios_cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket          (nios_cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready                (nios_cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid                (rsp_xbar_mux_src_valid),                                                                  //        rp.valid
		.rp_data                 (rsp_xbar_mux_src_data),                                                                   //          .data
		.rp_channel              (rsp_xbar_mux_src_channel),                                                                //          .channel
		.rp_startofpacket        (rsp_xbar_mux_src_startofpacket),                                                          //          .startofpacket
		.rp_endofpacket          (rsp_xbar_mux_src_endofpacket),                                                            //          .endofpacket
		.rp_ready                (rsp_xbar_mux_src_ready),                                                                  //          .ready
		.av_response             (),                                                                                        // (terminated)
		.av_writeresponserequest (1'b0),                                                                                    // (terminated)
		.av_writeresponsevalid   ()                                                                                         // (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_BEGIN_BURST           (77),
		.PKT_BURSTWRAP_H           (69),
		.PKT_BURSTWRAP_L           (67),
		.PKT_BURST_SIZE_H          (72),
		.PKT_BURST_SIZE_L          (70),
		.PKT_BURST_TYPE_H          (74),
		.PKT_BURST_TYPE_L          (73),
		.PKT_BYTE_CNT_H            (66),
		.PKT_BYTE_CNT_L            (64),
		.PKT_ADDR_H                (57),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (58),
		.PKT_TRANS_POSTED          (59),
		.PKT_TRANS_WRITE           (60),
		.PKT_TRANS_READ            (61),
		.PKT_TRANS_LOCK            (62),
		.PKT_TRANS_EXCLUSIVE       (63),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (85),
		.PKT_SRC_ID_L              (79),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (86),
		.PKT_THREAD_ID_H           (93),
		.PKT_THREAD_ID_L           (93),
		.PKT_CACHE_H               (100),
		.PKT_CACHE_L               (97),
		.PKT_DATA_SIDEBAND_H       (76),
		.PKT_DATA_SIDEBAND_L       (76),
		.PKT_QOS_H                 (78),
		.PKT_QOS_L                 (78),
		.PKT_ADDR_SIDEBAND_H       (75),
		.PKT_ADDR_SIDEBAND_L       (75),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.ST_DATA_W                 (103),
		.ST_CHANNEL_W              (99),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (0),
		.BURSTWRAP_VALUE           (7),
		.CACHE_VALUE               (0),
		.SECURE_ACCESS_BIT         (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) nios_cpu_data_master_translator_avalon_universal_master_0_agent (
		.clk                     (clk_clk),                                                                          //       clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                   // clk_reset.reset
		.av_address              (nios_cpu_data_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write                (nios_cpu_data_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read                 (nios_cpu_data_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata            (nios_cpu_data_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata             (nios_cpu_data_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest          (nios_cpu_data_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid        (nios_cpu_data_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable           (nios_cpu_data_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount           (nios_cpu_data_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess          (nios_cpu_data_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock                 (nios_cpu_data_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid                (nios_cpu_data_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data                 (nios_cpu_data_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket        (nios_cpu_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket          (nios_cpu_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready                (nios_cpu_data_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid                (rsp_xbar_mux_001_src_valid),                                                       //        rp.valid
		.rp_data                 (rsp_xbar_mux_001_src_data),                                                        //          .data
		.rp_channel              (rsp_xbar_mux_001_src_channel),                                                     //          .channel
		.rp_startofpacket        (rsp_xbar_mux_001_src_startofpacket),                                               //          .startofpacket
		.rp_endofpacket          (rsp_xbar_mux_001_src_endofpacket),                                                 //          .endofpacket
		.rp_ready                (rsp_xbar_mux_001_src_ready),                                                       //          .ready
		.av_response             (),                                                                                 // (terminated)
		.av_writeresponserequest (1'b0),                                                                             // (terminated)
		.av_writeresponsevalid   ()                                                                                  // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (77),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (57),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (58),
		.PKT_TRANS_POSTED          (59),
		.PKT_TRANS_WRITE           (60),
		.PKT_TRANS_READ            (61),
		.PKT_TRANS_LOCK            (62),
		.PKT_SRC_ID_H              (85),
		.PKT_SRC_ID_L              (79),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (86),
		.PKT_BURSTWRAP_H           (69),
		.PKT_BURSTWRAP_L           (67),
		.PKT_BYTE_CNT_H            (66),
		.PKT_BYTE_CNT_L            (64),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (72),
		.PKT_BURST_SIZE_L          (70),
		.ST_CHANNEL_W              (99),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) nios_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                         //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                  //       clk_reset.reset
		.m0_address              (nios_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (nios_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (nios_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (nios_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (nios_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (nios_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (nios_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (nios_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (nios_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (nios_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (nios_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (nios_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (nios_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (nios_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (nios_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (nios_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_src_ready),                                                                          //              cp.ready
		.cp_valid                (cmd_xbar_mux_src_valid),                                                                          //                .valid
		.cp_data                 (cmd_xbar_mux_src_data),                                                                           //                .data
		.cp_startofpacket        (cmd_xbar_mux_src_startofpacket),                                                                  //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_src_endofpacket),                                                                    //                .endofpacket
		.cp_channel              (cmd_xbar_mux_src_channel),                                                                        //                .channel
		.rf_sink_ready           (nios_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (nios_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (nios_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (nios_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (nios_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (nios_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (nios_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (nios_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (nios_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (nios_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (nios_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (nios_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (nios_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (nios_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (nios_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (nios_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                           //     (terminated)
		.m0_writeresponserequest (),                                                                                                //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                             //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) nios_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                         //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                  // clk_reset.reset
		.in_data           (nios_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (nios_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (nios_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (nios_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (nios_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (nios_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (nios_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (nios_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (nios_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (nios_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                           // (terminated)
		.csr_read          (1'b0),                                                                                            // (terminated)
		.csr_write         (1'b0),                                                                                            // (terminated)
		.csr_readdata      (),                                                                                                // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                            // (terminated)
		.almost_full_data  (),                                                                                                // (terminated)
		.almost_empty_data (),                                                                                                // (terminated)
		.in_empty          (1'b0),                                                                                            // (terminated)
		.out_empty         (),                                                                                                // (terminated)
		.in_error          (1'b0),                                                                                            // (terminated)
		.out_error         (),                                                                                                // (terminated)
		.in_channel        (1'b0),                                                                                            // (terminated)
		.out_channel       ()                                                                                                 // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (77),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (57),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (58),
		.PKT_TRANS_POSTED          (59),
		.PKT_TRANS_WRITE           (60),
		.PKT_TRANS_READ            (61),
		.PKT_TRANS_LOCK            (62),
		.PKT_SRC_ID_H              (85),
		.PKT_SRC_ID_L              (79),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (86),
		.PKT_BURSTWRAP_H           (69),
		.PKT_BURSTWRAP_L           (67),
		.PKT_BYTE_CNT_H            (66),
		.PKT_BYTE_CNT_L            (64),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (72),
		.PKT_BURST_SIZE_L          (70),
		.ST_CHANNEL_W              (99),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) ram_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                     //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                          //       clk_reset.reset
		.m0_address              (ram_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ram_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ram_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ram_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ram_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ram_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ram_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ram_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ram_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ram_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ram_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ram_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ram_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ram_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ram_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ram_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_001_src_ready),                                                  //              cp.ready
		.cp_valid                (cmd_xbar_mux_001_src_valid),                                                  //                .valid
		.cp_data                 (cmd_xbar_mux_001_src_data),                                                   //                .data
		.cp_startofpacket        (cmd_xbar_mux_001_src_startofpacket),                                          //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_001_src_endofpacket),                                            //                .endofpacket
		.cp_channel              (cmd_xbar_mux_001_src_channel),                                                //                .channel
		.rf_sink_ready           (ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ram_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ram_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ram_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ram_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ram_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (ram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (ram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                       //     (terminated)
		.m0_writeresponserequest (),                                                                            //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                         //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                     //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                          // clk_reset.reset
		.in_data           (ram_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ram_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ram_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ram_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ram_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                       // (terminated)
		.csr_read          (1'b0),                                                                        // (terminated)
		.csr_write         (1'b0),                                                                        // (terminated)
		.csr_readdata      (),                                                                            // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                        // (terminated)
		.almost_full_data  (),                                                                            // (terminated)
		.almost_empty_data (),                                                                            // (terminated)
		.in_empty          (1'b0),                                                                        // (terminated)
		.out_empty         (),                                                                            // (terminated)
		.in_error          (1'b0),                                                                        // (terminated)
		.out_error         (),                                                                            // (terminated)
		.in_channel        (1'b0),                                                                        // (terminated)
		.out_channel       ()                                                                             // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (77),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (57),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (58),
		.PKT_TRANS_POSTED          (59),
		.PKT_TRANS_WRITE           (60),
		.PKT_TRANS_READ            (61),
		.PKT_TRANS_LOCK            (62),
		.PKT_SRC_ID_H              (85),
		.PKT_SRC_ID_L              (79),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (86),
		.PKT_BURSTWRAP_H           (69),
		.PKT_BURSTWRAP_L           (67),
		.PKT_BYTE_CNT_H            (66),
		.PKT_BYTE_CNT_L            (64),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (72),
		.PKT_BURST_SIZE_L          (70),
		.ST_CHANNEL_W              (99),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) ssram_uas_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                        //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                             //       clk_reset.reset
		.m0_address              (ssram_uas_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ssram_uas_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ssram_uas_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ssram_uas_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ssram_uas_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ssram_uas_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ssram_uas_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ssram_uas_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ssram_uas_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ssram_uas_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ssram_uas_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ssram_uas_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ssram_uas_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ssram_uas_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ssram_uas_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ssram_uas_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_002_src_ready),                                                     //              cp.ready
		.cp_valid                (cmd_xbar_mux_002_src_valid),                                                     //                .valid
		.cp_data                 (cmd_xbar_mux_002_src_data),                                                      //                .data
		.cp_startofpacket        (cmd_xbar_mux_002_src_startofpacket),                                             //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_002_src_endofpacket),                                               //                .endofpacket
		.cp_channel              (cmd_xbar_mux_002_src_channel),                                                   //                .channel
		.rf_sink_ready           (ssram_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ssram_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ssram_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ssram_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ssram_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ssram_uas_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ssram_uas_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ssram_uas_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ssram_uas_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ssram_uas_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ssram_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ssram_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (ssram_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (ssram_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ssram_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ssram_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                          //     (terminated)
		.m0_writeresponserequest (),                                                                               //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                            //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (6),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ssram_uas_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                        //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                             // clk_reset.reset
		.in_data           (ssram_uas_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ssram_uas_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ssram_uas_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ssram_uas_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ssram_uas_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ssram_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ssram_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ssram_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ssram_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ssram_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                          // (terminated)
		.csr_read          (1'b0),                                                                           // (terminated)
		.csr_write         (1'b0),                                                                           // (terminated)
		.csr_readdata      (),                                                                               // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                           // (terminated)
		.almost_full_data  (),                                                                               // (terminated)
		.almost_empty_data (),                                                                               // (terminated)
		.in_empty          (1'b0),                                                                           // (terminated)
		.out_empty         (),                                                                               // (terminated)
		.in_error          (1'b0),                                                                           // (terminated)
		.out_error         (),                                                                               // (terminated)
		.in_channel        (1'b0),                                                                           // (terminated)
		.out_channel       ()                                                                                // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (77),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (57),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (58),
		.PKT_TRANS_POSTED          (59),
		.PKT_TRANS_WRITE           (60),
		.PKT_TRANS_READ            (61),
		.PKT_TRANS_LOCK            (62),
		.PKT_SRC_ID_H              (85),
		.PKT_SRC_ID_L              (79),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (86),
		.PKT_BURSTWRAP_H           (69),
		.PKT_BURSTWRAP_L           (67),
		.PKT_BYTE_CNT_H            (66),
		.PKT_BYTE_CNT_L            (64),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (72),
		.PKT_BURST_SIZE_L          (70),
		.ST_CHANNEL_W              (99),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                          //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                               //       clk_reset.reset
		.m0_address              (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src3_ready),                                                                    //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src3_valid),                                                                    //                .valid
		.cp_data                 (cmd_xbar_demux_001_src3_data),                                                                     //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src3_startofpacket),                                                            //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src3_endofpacket),                                                              //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src3_channel),                                                                  //                .channel
		.rf_sink_ready           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                            //     (terminated)
		.m0_writeresponserequest (),                                                                                                 //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                              //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                          //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                               // clk_reset.reset
		.in_data           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                            // (terminated)
		.csr_read          (1'b0),                                                                                             // (terminated)
		.csr_write         (1'b0),                                                                                             // (terminated)
		.csr_readdata      (),                                                                                                 // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                             // (terminated)
		.almost_full_data  (),                                                                                                 // (terminated)
		.almost_empty_data (),                                                                                                 // (terminated)
		.in_empty          (1'b0),                                                                                             // (terminated)
		.out_empty         (),                                                                                                 // (terminated)
		.in_error          (1'b0),                                                                                             // (terminated)
		.out_error         (),                                                                                                 // (terminated)
		.in_channel        (1'b0),                                                                                             // (terminated)
		.out_channel       ()                                                                                                  // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (77),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (57),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (58),
		.PKT_TRANS_POSTED          (59),
		.PKT_TRANS_WRITE           (60),
		.PKT_TRANS_READ            (61),
		.PKT_TRANS_LOCK            (62),
		.PKT_SRC_ID_H              (85),
		.PKT_SRC_ID_L              (79),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (86),
		.PKT_BURSTWRAP_H           (69),
		.PKT_BURSTWRAP_L           (67),
		.PKT_BYTE_CNT_H            (66),
		.PKT_BYTE_CNT_L            (64),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (72),
		.PKT_BURST_SIZE_L          (70),
		.ST_CHANNEL_W              (99),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) lcd_control_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                     //       clk_reset.reset
		.m0_address              (lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (lcd_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (lcd_control_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (lcd_control_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (lcd_control_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (lcd_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src4_ready),                                                          //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src4_valid),                                                          //                .valid
		.cp_data                 (cmd_xbar_demux_001_src4_data),                                                           //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src4_startofpacket),                                                  //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src4_endofpacket),                                                    //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src4_channel),                                                        //                .channel
		.rf_sink_ready           (lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (lcd_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (lcd_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (lcd_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (lcd_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (lcd_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (lcd_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (lcd_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (lcd_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (lcd_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (lcd_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (lcd_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                  //     (terminated)
		.m0_writeresponserequest (),                                                                                       //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                    //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                     // clk_reset.reset
		.in_data           (lcd_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (lcd_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (lcd_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (lcd_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (lcd_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                  // (terminated)
		.csr_read          (1'b0),                                                                                   // (terminated)
		.csr_write         (1'b0),                                                                                   // (terminated)
		.csr_readdata      (),                                                                                       // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                   // (terminated)
		.almost_full_data  (),                                                                                       // (terminated)
		.almost_empty_data (),                                                                                       // (terminated)
		.in_empty          (1'b0),                                                                                   // (terminated)
		.out_empty         (),                                                                                       // (terminated)
		.in_error          (1'b0),                                                                                   // (terminated)
		.out_error         (),                                                                                       // (terminated)
		.in_channel        (1'b0),                                                                                   // (terminated)
		.out_channel       ()                                                                                        // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (77),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (57),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (58),
		.PKT_TRANS_POSTED          (59),
		.PKT_TRANS_WRITE           (60),
		.PKT_TRANS_READ            (61),
		.PKT_TRANS_LOCK            (62),
		.PKT_SRC_ID_H              (85),
		.PKT_SRC_ID_L              (79),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (86),
		.PKT_BURSTWRAP_H           (69),
		.PKT_BURSTWRAP_L           (67),
		.PKT_BYTE_CNT_H            (66),
		.PKT_BYTE_CNT_L            (64),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (72),
		.PKT_BURST_SIZE_L          (70),
		.ST_CHANNEL_W              (99),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) adc_on_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                        //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                             //       clk_reset.reset
		.m0_address              (adc_on_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (adc_on_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (adc_on_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (adc_on_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (adc_on_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (adc_on_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (adc_on_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (adc_on_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (adc_on_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (adc_on_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (adc_on_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (adc_on_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (adc_on_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (adc_on_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (adc_on_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (adc_on_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src5_ready),                                                  //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src5_valid),                                                  //                .valid
		.cp_data                 (cmd_xbar_demux_001_src5_data),                                                   //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src5_startofpacket),                                          //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src5_endofpacket),                                            //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src5_channel),                                                //                .channel
		.rf_sink_ready           (adc_on_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (adc_on_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (adc_on_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (adc_on_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (adc_on_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (adc_on_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (adc_on_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (adc_on_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (adc_on_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (adc_on_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (adc_on_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (adc_on_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (adc_on_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (adc_on_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (adc_on_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (adc_on_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                          //     (terminated)
		.m0_writeresponserequest (),                                                                               //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                            //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) adc_on_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                        //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                             // clk_reset.reset
		.in_data           (adc_on_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (adc_on_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (adc_on_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (adc_on_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (adc_on_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (adc_on_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (adc_on_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (adc_on_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (adc_on_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (adc_on_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                          // (terminated)
		.csr_read          (1'b0),                                                                           // (terminated)
		.csr_write         (1'b0),                                                                           // (terminated)
		.csr_readdata      (),                                                                               // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                           // (terminated)
		.almost_full_data  (),                                                                               // (terminated)
		.almost_empty_data (),                                                                               // (terminated)
		.in_empty          (1'b0),                                                                           // (terminated)
		.out_empty         (),                                                                               // (terminated)
		.in_error          (1'b0),                                                                           // (terminated)
		.out_error         (),                                                                               // (terminated)
		.in_channel        (1'b0),                                                                           // (terminated)
		.out_channel       ()                                                                                // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (77),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (57),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (58),
		.PKT_TRANS_POSTED          (59),
		.PKT_TRANS_WRITE           (60),
		.PKT_TRANS_READ            (61),
		.PKT_TRANS_LOCK            (62),
		.PKT_SRC_ID_H              (85),
		.PKT_SRC_ID_L              (79),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (86),
		.PKT_BURSTWRAP_H           (69),
		.PKT_BURSTWRAP_L           (67),
		.PKT_BYTE_CNT_H            (66),
		.PKT_BYTE_CNT_L            (64),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (72),
		.PKT_BURST_SIZE_L          (70),
		.ST_CHANNEL_W              (99),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) fifo_adc_data_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                               //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                    //       clk_reset.reset
		.m0_address              (fifo_adc_data_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (fifo_adc_data_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (fifo_adc_data_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (fifo_adc_data_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (fifo_adc_data_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (fifo_adc_data_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (fifo_adc_data_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (fifo_adc_data_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (fifo_adc_data_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (fifo_adc_data_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (fifo_adc_data_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (fifo_adc_data_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (fifo_adc_data_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (fifo_adc_data_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (fifo_adc_data_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (fifo_adc_data_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src6_ready),                                                         //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src6_valid),                                                         //                .valid
		.cp_data                 (cmd_xbar_demux_001_src6_data),                                                          //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src6_startofpacket),                                                 //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src6_endofpacket),                                                   //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src6_channel),                                                       //                .channel
		.rf_sink_ready           (fifo_adc_data_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (fifo_adc_data_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (fifo_adc_data_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (fifo_adc_data_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (fifo_adc_data_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (fifo_adc_data_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (fifo_adc_data_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (fifo_adc_data_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (fifo_adc_data_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (fifo_adc_data_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (fifo_adc_data_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (fifo_adc_data_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (fifo_adc_data_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (fifo_adc_data_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (fifo_adc_data_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (fifo_adc_data_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                 //     (terminated)
		.m0_writeresponserequest (),                                                                                      //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                   //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) fifo_adc_data_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                               //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                    // clk_reset.reset
		.in_data           (fifo_adc_data_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (fifo_adc_data_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (fifo_adc_data_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (fifo_adc_data_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (fifo_adc_data_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (fifo_adc_data_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (fifo_adc_data_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (fifo_adc_data_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (fifo_adc_data_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (fifo_adc_data_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                 // (terminated)
		.csr_read          (1'b0),                                                                                  // (terminated)
		.csr_write         (1'b0),                                                                                  // (terminated)
		.csr_readdata      (),                                                                                      // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                  // (terminated)
		.almost_full_data  (),                                                                                      // (terminated)
		.almost_empty_data (),                                                                                      // (terminated)
		.in_empty          (1'b0),                                                                                  // (terminated)
		.out_empty         (),                                                                                      // (terminated)
		.in_error          (1'b0),                                                                                  // (terminated)
		.out_error         (),                                                                                      // (terminated)
		.in_channel        (1'b0),                                                                                  // (terminated)
		.out_channel       ()                                                                                       // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (77),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (57),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (58),
		.PKT_TRANS_POSTED          (59),
		.PKT_TRANS_WRITE           (60),
		.PKT_TRANS_READ            (61),
		.PKT_TRANS_LOCK            (62),
		.PKT_SRC_ID_H              (85),
		.PKT_SRC_ID_L              (79),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (86),
		.PKT_BURSTWRAP_H           (69),
		.PKT_BURSTWRAP_L           (67),
		.PKT_BYTE_CNT_H            (66),
		.PKT_BYTE_CNT_L            (64),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (72),
		.PKT_BURST_SIZE_L          (70),
		.ST_CHANNEL_W              (99),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) fifo_adc_data_valid_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                     //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                          //       clk_reset.reset
		.m0_address              (fifo_adc_data_valid_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (fifo_adc_data_valid_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (fifo_adc_data_valid_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (fifo_adc_data_valid_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (fifo_adc_data_valid_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (fifo_adc_data_valid_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (fifo_adc_data_valid_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (fifo_adc_data_valid_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (fifo_adc_data_valid_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (fifo_adc_data_valid_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (fifo_adc_data_valid_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (fifo_adc_data_valid_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (fifo_adc_data_valid_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (fifo_adc_data_valid_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (fifo_adc_data_valid_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (fifo_adc_data_valid_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src7_ready),                                                               //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src7_valid),                                                               //                .valid
		.cp_data                 (cmd_xbar_demux_001_src7_data),                                                                //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src7_startofpacket),                                                       //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src7_endofpacket),                                                         //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src7_channel),                                                             //                .channel
		.rf_sink_ready           (fifo_adc_data_valid_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (fifo_adc_data_valid_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (fifo_adc_data_valid_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (fifo_adc_data_valid_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (fifo_adc_data_valid_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (fifo_adc_data_valid_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (fifo_adc_data_valid_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (fifo_adc_data_valid_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (fifo_adc_data_valid_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (fifo_adc_data_valid_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (fifo_adc_data_valid_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (fifo_adc_data_valid_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (fifo_adc_data_valid_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (fifo_adc_data_valid_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (fifo_adc_data_valid_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (fifo_adc_data_valid_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                       //     (terminated)
		.m0_writeresponserequest (),                                                                                            //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                         //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) fifo_adc_data_valid_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                     //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                          // clk_reset.reset
		.in_data           (fifo_adc_data_valid_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (fifo_adc_data_valid_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (fifo_adc_data_valid_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (fifo_adc_data_valid_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (fifo_adc_data_valid_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (fifo_adc_data_valid_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (fifo_adc_data_valid_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (fifo_adc_data_valid_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (fifo_adc_data_valid_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (fifo_adc_data_valid_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                       // (terminated)
		.csr_read          (1'b0),                                                                                        // (terminated)
		.csr_write         (1'b0),                                                                                        // (terminated)
		.csr_readdata      (),                                                                                            // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                        // (terminated)
		.almost_full_data  (),                                                                                            // (terminated)
		.almost_empty_data (),                                                                                            // (terminated)
		.in_empty          (1'b0),                                                                                        // (terminated)
		.out_empty         (),                                                                                            // (terminated)
		.in_error          (1'b0),                                                                                        // (terminated)
		.out_error         (),                                                                                            // (terminated)
		.in_channel        (1'b0),                                                                                        // (terminated)
		.out_channel       ()                                                                                             // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (77),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (57),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (58),
		.PKT_TRANS_POSTED          (59),
		.PKT_TRANS_WRITE           (60),
		.PKT_TRANS_READ            (61),
		.PKT_TRANS_LOCK            (62),
		.PKT_SRC_ID_H              (85),
		.PKT_SRC_ID_L              (79),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (86),
		.PKT_BURSTWRAP_H           (69),
		.PKT_BURSTWRAP_L           (67),
		.PKT_BYTE_CNT_H            (66),
		.PKT_BYTE_CNT_L            (64),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (72),
		.PKT_BURST_SIZE_L          (70),
		.ST_CHANNEL_W              (99),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) fifo_rst_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                          //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                               //       clk_reset.reset
		.m0_address              (fifo_rst_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (fifo_rst_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (fifo_rst_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (fifo_rst_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (fifo_rst_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (fifo_rst_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (fifo_rst_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (fifo_rst_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (fifo_rst_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (fifo_rst_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (fifo_rst_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (fifo_rst_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (fifo_rst_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (fifo_rst_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (fifo_rst_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (fifo_rst_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src8_ready),                                                    //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src8_valid),                                                    //                .valid
		.cp_data                 (cmd_xbar_demux_001_src8_data),                                                     //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src8_startofpacket),                                            //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src8_endofpacket),                                              //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src8_channel),                                                  //                .channel
		.rf_sink_ready           (fifo_rst_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (fifo_rst_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (fifo_rst_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (fifo_rst_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (fifo_rst_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (fifo_rst_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (fifo_rst_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (fifo_rst_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (fifo_rst_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (fifo_rst_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (fifo_rst_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (fifo_rst_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (fifo_rst_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (fifo_rst_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (fifo_rst_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (fifo_rst_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                            //     (terminated)
		.m0_writeresponserequest (),                                                                                 //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                              //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) fifo_rst_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                          //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                               // clk_reset.reset
		.in_data           (fifo_rst_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (fifo_rst_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (fifo_rst_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (fifo_rst_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (fifo_rst_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (fifo_rst_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (fifo_rst_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (fifo_rst_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (fifo_rst_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (fifo_rst_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                            // (terminated)
		.csr_read          (1'b0),                                                                             // (terminated)
		.csr_write         (1'b0),                                                                             // (terminated)
		.csr_readdata      (),                                                                                 // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                             // (terminated)
		.almost_full_data  (),                                                                                 // (terminated)
		.almost_empty_data (),                                                                                 // (terminated)
		.in_empty          (1'b0),                                                                             // (terminated)
		.out_empty         (),                                                                                 // (terminated)
		.in_error          (1'b0),                                                                             // (terminated)
		.out_error         (),                                                                                 // (terminated)
		.in_channel        (1'b0),                                                                             // (terminated)
		.out_channel       ()                                                                                  // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (77),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (57),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (58),
		.PKT_TRANS_POSTED          (59),
		.PKT_TRANS_WRITE           (60),
		.PKT_TRANS_READ            (61),
		.PKT_TRANS_LOCK            (62),
		.PKT_SRC_ID_H              (85),
		.PKT_SRC_ID_L              (79),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (86),
		.PKT_BURSTWRAP_H           (69),
		.PKT_BURSTWRAP_L           (67),
		.PKT_BYTE_CNT_H            (66),
		.PKT_BYTE_CNT_L            (64),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (72),
		.PKT_BURST_SIZE_L          (70),
		.ST_CHANNEL_W              (99),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) subtractor_on_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                               //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                    //       clk_reset.reset
		.m0_address              (subtractor_on_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (subtractor_on_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (subtractor_on_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (subtractor_on_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (subtractor_on_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (subtractor_on_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (subtractor_on_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (subtractor_on_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (subtractor_on_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (subtractor_on_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (subtractor_on_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (subtractor_on_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (subtractor_on_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (subtractor_on_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (subtractor_on_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (subtractor_on_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src9_ready),                                                         //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src9_valid),                                                         //                .valid
		.cp_data                 (cmd_xbar_demux_001_src9_data),                                                          //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src9_startofpacket),                                                 //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src9_endofpacket),                                                   //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src9_channel),                                                       //                .channel
		.rf_sink_ready           (subtractor_on_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (subtractor_on_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (subtractor_on_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (subtractor_on_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (subtractor_on_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (subtractor_on_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (subtractor_on_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (subtractor_on_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (subtractor_on_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (subtractor_on_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (subtractor_on_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (subtractor_on_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (subtractor_on_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (subtractor_on_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (subtractor_on_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (subtractor_on_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                 //     (terminated)
		.m0_writeresponserequest (),                                                                                      //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                   //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) subtractor_on_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                               //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                    // clk_reset.reset
		.in_data           (subtractor_on_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (subtractor_on_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (subtractor_on_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (subtractor_on_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (subtractor_on_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (subtractor_on_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (subtractor_on_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (subtractor_on_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (subtractor_on_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (subtractor_on_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                 // (terminated)
		.csr_read          (1'b0),                                                                                  // (terminated)
		.csr_write         (1'b0),                                                                                  // (terminated)
		.csr_readdata      (),                                                                                      // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                  // (terminated)
		.almost_full_data  (),                                                                                      // (terminated)
		.almost_empty_data (),                                                                                      // (terminated)
		.in_empty          (1'b0),                                                                                  // (terminated)
		.out_empty         (),                                                                                      // (terminated)
		.in_error          (1'b0),                                                                                  // (terminated)
		.out_error         (),                                                                                      // (terminated)
		.in_channel        (1'b0),                                                                                  // (terminated)
		.out_channel       ()                                                                                       // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (77),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (57),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (58),
		.PKT_TRANS_POSTED          (59),
		.PKT_TRANS_WRITE           (60),
		.PKT_TRANS_READ            (61),
		.PKT_TRANS_LOCK            (62),
		.PKT_SRC_ID_H              (85),
		.PKT_SRC_ID_L              (79),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (86),
		.PKT_BURSTWRAP_H           (69),
		.PKT_BURSTWRAP_L           (67),
		.PKT_BYTE_CNT_H            (66),
		.PKT_BYTE_CNT_L            (64),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (72),
		.PKT_BURST_SIZE_L          (70),
		.ST_CHANNEL_W              (99),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) ch0_timer_rst_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                               //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                    //       clk_reset.reset
		.m0_address              (ch0_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ch0_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ch0_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ch0_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ch0_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ch0_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ch0_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ch0_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ch0_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ch0_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ch0_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ch0_timer_rst_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ch0_timer_rst_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ch0_timer_rst_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ch0_timer_rst_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ch0_timer_rst_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src10_ready),                                                        //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src10_valid),                                                        //                .valid
		.cp_data                 (cmd_xbar_demux_001_src10_data),                                                         //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src10_startofpacket),                                                //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src10_endofpacket),                                                  //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src10_channel),                                                      //                .channel
		.rf_sink_ready           (ch0_timer_rst_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ch0_timer_rst_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ch0_timer_rst_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ch0_timer_rst_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ch0_timer_rst_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ch0_timer_rst_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ch0_timer_rst_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ch0_timer_rst_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ch0_timer_rst_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ch0_timer_rst_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ch0_timer_rst_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ch0_timer_rst_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (ch0_timer_rst_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (ch0_timer_rst_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ch0_timer_rst_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ch0_timer_rst_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                 //     (terminated)
		.m0_writeresponserequest (),                                                                                      //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                   //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ch0_timer_rst_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                               //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                    // clk_reset.reset
		.in_data           (ch0_timer_rst_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ch0_timer_rst_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ch0_timer_rst_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ch0_timer_rst_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ch0_timer_rst_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ch0_timer_rst_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ch0_timer_rst_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ch0_timer_rst_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ch0_timer_rst_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ch0_timer_rst_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                 // (terminated)
		.csr_read          (1'b0),                                                                                  // (terminated)
		.csr_write         (1'b0),                                                                                  // (terminated)
		.csr_readdata      (),                                                                                      // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                  // (terminated)
		.almost_full_data  (),                                                                                      // (terminated)
		.almost_empty_data (),                                                                                      // (terminated)
		.in_empty          (1'b0),                                                                                  // (terminated)
		.out_empty         (),                                                                                      // (terminated)
		.in_error          (1'b0),                                                                                  // (terminated)
		.out_error         (),                                                                                      // (terminated)
		.in_channel        (1'b0),                                                                                  // (terminated)
		.out_channel       ()                                                                                       // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (77),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (57),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (58),
		.PKT_TRANS_POSTED          (59),
		.PKT_TRANS_WRITE           (60),
		.PKT_TRANS_READ            (61),
		.PKT_TRANS_LOCK            (62),
		.PKT_SRC_ID_H              (85),
		.PKT_SRC_ID_L              (79),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (86),
		.PKT_BURSTWRAP_H           (69),
		.PKT_BURSTWRAP_L           (67),
		.PKT_BYTE_CNT_H            (66),
		.PKT_BYTE_CNT_L            (64),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (72),
		.PKT_BURST_SIZE_L          (70),
		.ST_CHANNEL_W              (99),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) detector_on_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                             //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                  //       clk_reset.reset
		.m0_address              (detector_on_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (detector_on_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (detector_on_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (detector_on_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (detector_on_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (detector_on_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (detector_on_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (detector_on_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (detector_on_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (detector_on_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (detector_on_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (detector_on_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (detector_on_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (detector_on_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (detector_on_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (detector_on_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src11_ready),                                                      //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src11_valid),                                                      //                .valid
		.cp_data                 (cmd_xbar_demux_001_src11_data),                                                       //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src11_startofpacket),                                              //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src11_endofpacket),                                                //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src11_channel),                                                    //                .channel
		.rf_sink_ready           (detector_on_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (detector_on_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (detector_on_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (detector_on_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (detector_on_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (detector_on_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (detector_on_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (detector_on_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (detector_on_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (detector_on_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (detector_on_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (detector_on_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (detector_on_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (detector_on_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (detector_on_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (detector_on_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                               //     (terminated)
		.m0_writeresponserequest (),                                                                                    //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                 //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) detector_on_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                             //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                  // clk_reset.reset
		.in_data           (detector_on_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (detector_on_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (detector_on_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (detector_on_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (detector_on_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (detector_on_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (detector_on_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (detector_on_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (detector_on_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (detector_on_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                               // (terminated)
		.csr_read          (1'b0),                                                                                // (terminated)
		.csr_write         (1'b0),                                                                                // (terminated)
		.csr_readdata      (),                                                                                    // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                // (terminated)
		.almost_full_data  (),                                                                                    // (terminated)
		.almost_empty_data (),                                                                                    // (terminated)
		.in_empty          (1'b0),                                                                                // (terminated)
		.out_empty         (),                                                                                    // (terminated)
		.in_error          (1'b0),                                                                                // (terminated)
		.out_error         (),                                                                                    // (terminated)
		.in_channel        (1'b0),                                                                                // (terminated)
		.out_channel       ()                                                                                     // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (77),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (57),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (58),
		.PKT_TRANS_POSTED          (59),
		.PKT_TRANS_WRITE           (60),
		.PKT_TRANS_READ            (61),
		.PKT_TRANS_LOCK            (62),
		.PKT_SRC_ID_H              (85),
		.PKT_SRC_ID_L              (79),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (86),
		.PKT_BURSTWRAP_H           (69),
		.PKT_BURSTWRAP_L           (67),
		.PKT_BYTE_CNT_H            (66),
		.PKT_BYTE_CNT_L            (64),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (72),
		.PKT_BURST_SIZE_L          (70),
		.ST_CHANNEL_W              (99),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) menu_down_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                           //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                //       clk_reset.reset
		.m0_address              (menu_down_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (menu_down_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (menu_down_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (menu_down_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (menu_down_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (menu_down_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (menu_down_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (menu_down_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (menu_down_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (menu_down_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (menu_down_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (menu_down_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (menu_down_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (menu_down_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (menu_down_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (menu_down_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src12_ready),                                                    //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src12_valid),                                                    //                .valid
		.cp_data                 (cmd_xbar_demux_001_src12_data),                                                     //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src12_startofpacket),                                            //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src12_endofpacket),                                              //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src12_channel),                                                  //                .channel
		.rf_sink_ready           (menu_down_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (menu_down_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (menu_down_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (menu_down_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (menu_down_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (menu_down_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (menu_down_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (menu_down_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (menu_down_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (menu_down_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (menu_down_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (menu_down_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (menu_down_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (menu_down_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (menu_down_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (menu_down_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                             //     (terminated)
		.m0_writeresponserequest (),                                                                                  //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                               //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) menu_down_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                           //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                // clk_reset.reset
		.in_data           (menu_down_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (menu_down_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (menu_down_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (menu_down_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (menu_down_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (menu_down_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (menu_down_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (menu_down_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (menu_down_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (menu_down_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                             // (terminated)
		.csr_read          (1'b0),                                                                              // (terminated)
		.csr_write         (1'b0),                                                                              // (terminated)
		.csr_readdata      (),                                                                                  // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                              // (terminated)
		.almost_full_data  (),                                                                                  // (terminated)
		.almost_empty_data (),                                                                                  // (terminated)
		.in_empty          (1'b0),                                                                              // (terminated)
		.out_empty         (),                                                                                  // (terminated)
		.in_error          (1'b0),                                                                              // (terminated)
		.out_error         (),                                                                                  // (terminated)
		.in_channel        (1'b0),                                                                              // (terminated)
		.out_channel       ()                                                                                   // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (77),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (57),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (58),
		.PKT_TRANS_POSTED          (59),
		.PKT_TRANS_WRITE           (60),
		.PKT_TRANS_READ            (61),
		.PKT_TRANS_LOCK            (62),
		.PKT_SRC_ID_H              (85),
		.PKT_SRC_ID_L              (79),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (86),
		.PKT_BURSTWRAP_H           (69),
		.PKT_BURSTWRAP_L           (67),
		.PKT_BYTE_CNT_H            (66),
		.PKT_BYTE_CNT_L            (64),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (72),
		.PKT_BURST_SIZE_L          (70),
		.ST_CHANNEL_W              (99),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) menu_up_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                         //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                              //       clk_reset.reset
		.m0_address              (menu_up_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (menu_up_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (menu_up_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (menu_up_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (menu_up_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (menu_up_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (menu_up_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (menu_up_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (menu_up_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (menu_up_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (menu_up_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (menu_up_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (menu_up_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (menu_up_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (menu_up_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (menu_up_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src13_ready),                                                  //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src13_valid),                                                  //                .valid
		.cp_data                 (cmd_xbar_demux_001_src13_data),                                                   //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src13_startofpacket),                                          //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src13_endofpacket),                                            //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src13_channel),                                                //                .channel
		.rf_sink_ready           (menu_up_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (menu_up_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (menu_up_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (menu_up_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (menu_up_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (menu_up_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (menu_up_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (menu_up_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (menu_up_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (menu_up_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (menu_up_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (menu_up_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (menu_up_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (menu_up_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (menu_up_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (menu_up_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                           //     (terminated)
		.m0_writeresponserequest (),                                                                                //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                             //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) menu_up_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                         //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                              // clk_reset.reset
		.in_data           (menu_up_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (menu_up_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (menu_up_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (menu_up_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (menu_up_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (menu_up_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (menu_up_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (menu_up_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (menu_up_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (menu_up_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                           // (terminated)
		.csr_read          (1'b0),                                                                            // (terminated)
		.csr_write         (1'b0),                                                                            // (terminated)
		.csr_readdata      (),                                                                                // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                            // (terminated)
		.almost_full_data  (),                                                                                // (terminated)
		.almost_empty_data (),                                                                                // (terminated)
		.in_empty          (1'b0),                                                                            // (terminated)
		.out_empty         (),                                                                                // (terminated)
		.in_error          (1'b0),                                                                            // (terminated)
		.out_error         (),                                                                                // (terminated)
		.in_channel        (1'b0),                                                                            // (terminated)
		.out_channel       ()                                                                                 // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (77),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (57),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (58),
		.PKT_TRANS_POSTED          (59),
		.PKT_TRANS_WRITE           (60),
		.PKT_TRANS_READ            (61),
		.PKT_TRANS_LOCK            (62),
		.PKT_SRC_ID_H              (85),
		.PKT_SRC_ID_L              (79),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (86),
		.PKT_BURSTWRAP_H           (69),
		.PKT_BURSTWRAP_L           (67),
		.PKT_BYTE_CNT_H            (66),
		.PKT_BYTE_CNT_L            (64),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (72),
		.PKT_BURST_SIZE_L          (70),
		.ST_CHANNEL_W              (99),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) menu_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                      //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                           //       clk_reset.reset
		.m0_address              (menu_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (menu_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (menu_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (menu_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (menu_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (menu_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (menu_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (menu_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (menu_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (menu_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (menu_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (menu_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (menu_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (menu_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (menu_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (menu_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src14_ready),                                               //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src14_valid),                                               //                .valid
		.cp_data                 (cmd_xbar_demux_001_src14_data),                                                //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src14_startofpacket),                                       //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src14_endofpacket),                                         //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src14_channel),                                             //                .channel
		.rf_sink_ready           (menu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (menu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (menu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (menu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (menu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (menu_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (menu_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (menu_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (menu_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (menu_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (menu_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (menu_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (menu_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (menu_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (menu_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (menu_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                        //     (terminated)
		.m0_writeresponserequest (),                                                                             //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                          //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) menu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                      //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                           // clk_reset.reset
		.in_data           (menu_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (menu_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (menu_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (menu_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (menu_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (menu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (menu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (menu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (menu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (menu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                        // (terminated)
		.csr_read          (1'b0),                                                                         // (terminated)
		.csr_write         (1'b0),                                                                         // (terminated)
		.csr_readdata      (),                                                                             // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                         // (terminated)
		.almost_full_data  (),                                                                             // (terminated)
		.almost_empty_data (),                                                                             // (terminated)
		.in_empty          (1'b0),                                                                         // (terminated)
		.out_empty         (),                                                                             // (terminated)
		.in_error          (1'b0),                                                                         // (terminated)
		.out_error         (),                                                                             // (terminated)
		.in_channel        (1'b0),                                                                         // (terminated)
		.out_channel       ()                                                                              // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (77),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (57),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (58),
		.PKT_TRANS_POSTED          (59),
		.PKT_TRANS_WRITE           (60),
		.PKT_TRANS_READ            (61),
		.PKT_TRANS_LOCK            (62),
		.PKT_SRC_ID_H              (85),
		.PKT_SRC_ID_L              (79),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (86),
		.PKT_BURSTWRAP_H           (69),
		.PKT_BURSTWRAP_L           (67),
		.PKT_BYTE_CNT_H            (66),
		.PKT_BYTE_CNT_L            (64),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (72),
		.PKT_BURST_SIZE_L          (70),
		.ST_CHANNEL_W              (99),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) ch0_thresh_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                            //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                 //       clk_reset.reset
		.m0_address              (ch0_thresh_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ch0_thresh_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ch0_thresh_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ch0_thresh_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ch0_thresh_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ch0_thresh_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ch0_thresh_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ch0_thresh_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ch0_thresh_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ch0_thresh_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ch0_thresh_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ch0_thresh_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ch0_thresh_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ch0_thresh_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ch0_thresh_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ch0_thresh_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src15_ready),                                                     //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src15_valid),                                                     //                .valid
		.cp_data                 (cmd_xbar_demux_001_src15_data),                                                      //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src15_startofpacket),                                             //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src15_endofpacket),                                               //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src15_channel),                                                   //                .channel
		.rf_sink_ready           (ch0_thresh_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ch0_thresh_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ch0_thresh_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ch0_thresh_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ch0_thresh_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ch0_thresh_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ch0_thresh_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ch0_thresh_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ch0_thresh_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ch0_thresh_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ch0_thresh_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ch0_thresh_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (ch0_thresh_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (ch0_thresh_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ch0_thresh_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ch0_thresh_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                              //     (terminated)
		.m0_writeresponserequest (),                                                                                   //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ch0_thresh_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                            //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                 // clk_reset.reset
		.in_data           (ch0_thresh_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ch0_thresh_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ch0_thresh_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ch0_thresh_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ch0_thresh_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ch0_thresh_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ch0_thresh_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ch0_thresh_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ch0_thresh_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ch0_thresh_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                              // (terminated)
		.csr_read          (1'b0),                                                                               // (terminated)
		.csr_write         (1'b0),                                                                               // (terminated)
		.csr_readdata      (),                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                               // (terminated)
		.almost_full_data  (),                                                                                   // (terminated)
		.almost_empty_data (),                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                               // (terminated)
		.out_empty         (),                                                                                   // (terminated)
		.in_error          (1'b0),                                                                               // (terminated)
		.out_error         (),                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                               // (terminated)
		.out_channel       ()                                                                                    // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (77),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (57),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (58),
		.PKT_TRANS_POSTED          (59),
		.PKT_TRANS_WRITE           (60),
		.PKT_TRANS_READ            (61),
		.PKT_TRANS_LOCK            (62),
		.PKT_SRC_ID_H              (85),
		.PKT_SRC_ID_L              (79),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (86),
		.PKT_BURSTWRAP_H           (69),
		.PKT_BURSTWRAP_L           (67),
		.PKT_BYTE_CNT_H            (66),
		.PKT_BYTE_CNT_L            (64),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (72),
		.PKT_BURST_SIZE_L          (70),
		.ST_CHANNEL_W              (99),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) ch0_rd_peak_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                             //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                  //       clk_reset.reset
		.m0_address              (ch0_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ch0_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ch0_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ch0_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ch0_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ch0_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ch0_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ch0_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ch0_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ch0_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ch0_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ch0_rd_peak_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ch0_rd_peak_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ch0_rd_peak_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ch0_rd_peak_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ch0_rd_peak_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src16_ready),                                                      //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src16_valid),                                                      //                .valid
		.cp_data                 (cmd_xbar_demux_001_src16_data),                                                       //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src16_startofpacket),                                              //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src16_endofpacket),                                                //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src16_channel),                                                    //                .channel
		.rf_sink_ready           (ch0_rd_peak_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ch0_rd_peak_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ch0_rd_peak_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ch0_rd_peak_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ch0_rd_peak_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ch0_rd_peak_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ch0_rd_peak_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ch0_rd_peak_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ch0_rd_peak_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ch0_rd_peak_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ch0_rd_peak_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ch0_rd_peak_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (ch0_rd_peak_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (ch0_rd_peak_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ch0_rd_peak_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ch0_rd_peak_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                               //     (terminated)
		.m0_writeresponserequest (),                                                                                    //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                 //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ch0_rd_peak_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                             //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                  // clk_reset.reset
		.in_data           (ch0_rd_peak_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ch0_rd_peak_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ch0_rd_peak_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ch0_rd_peak_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ch0_rd_peak_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ch0_rd_peak_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ch0_rd_peak_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ch0_rd_peak_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ch0_rd_peak_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ch0_rd_peak_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                               // (terminated)
		.csr_read          (1'b0),                                                                                // (terminated)
		.csr_write         (1'b0),                                                                                // (terminated)
		.csr_readdata      (),                                                                                    // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                // (terminated)
		.almost_full_data  (),                                                                                    // (terminated)
		.almost_empty_data (),                                                                                    // (terminated)
		.in_empty          (1'b0),                                                                                // (terminated)
		.out_empty         (),                                                                                    // (terminated)
		.in_error          (1'b0),                                                                                // (terminated)
		.out_error         (),                                                                                    // (terminated)
		.in_channel        (1'b0),                                                                                // (terminated)
		.out_channel       ()                                                                                     // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (77),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (57),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (58),
		.PKT_TRANS_POSTED          (59),
		.PKT_TRANS_WRITE           (60),
		.PKT_TRANS_READ            (61),
		.PKT_TRANS_LOCK            (62),
		.PKT_SRC_ID_H              (85),
		.PKT_SRC_ID_L              (79),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (86),
		.PKT_BURSTWRAP_H           (69),
		.PKT_BURSTWRAP_L           (67),
		.PKT_BYTE_CNT_H            (66),
		.PKT_BYTE_CNT_L            (64),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (72),
		.PKT_BURST_SIZE_L          (70),
		.ST_CHANNEL_W              (99),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) ch0_peak_found_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                     //       clk_reset.reset
		.m0_address              (ch0_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ch0_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ch0_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ch0_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ch0_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ch0_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ch0_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ch0_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ch0_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ch0_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ch0_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ch0_peak_found_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ch0_peak_found_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ch0_peak_found_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ch0_peak_found_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ch0_peak_found_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src17_ready),                                                         //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src17_valid),                                                         //                .valid
		.cp_data                 (cmd_xbar_demux_001_src17_data),                                                          //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src17_startofpacket),                                                 //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src17_endofpacket),                                                   //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src17_channel),                                                       //                .channel
		.rf_sink_ready           (ch0_peak_found_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ch0_peak_found_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ch0_peak_found_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ch0_peak_found_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ch0_peak_found_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ch0_peak_found_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ch0_peak_found_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ch0_peak_found_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ch0_peak_found_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ch0_peak_found_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ch0_peak_found_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ch0_peak_found_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (ch0_peak_found_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (ch0_peak_found_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ch0_peak_found_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ch0_peak_found_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                  //     (terminated)
		.m0_writeresponserequest (),                                                                                       //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                    //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ch0_peak_found_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                     // clk_reset.reset
		.in_data           (ch0_peak_found_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ch0_peak_found_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ch0_peak_found_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ch0_peak_found_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ch0_peak_found_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ch0_peak_found_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ch0_peak_found_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ch0_peak_found_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ch0_peak_found_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ch0_peak_found_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                  // (terminated)
		.csr_read          (1'b0),                                                                                   // (terminated)
		.csr_write         (1'b0),                                                                                   // (terminated)
		.csr_readdata      (),                                                                                       // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                   // (terminated)
		.almost_full_data  (),                                                                                       // (terminated)
		.almost_empty_data (),                                                                                       // (terminated)
		.in_empty          (1'b0),                                                                                   // (terminated)
		.out_empty         (),                                                                                       // (terminated)
		.in_error          (1'b0),                                                                                   // (terminated)
		.out_error         (),                                                                                       // (terminated)
		.in_channel        (1'b0),                                                                                   // (terminated)
		.out_channel       ()                                                                                        // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (77),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (57),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (58),
		.PKT_TRANS_POSTED          (59),
		.PKT_TRANS_WRITE           (60),
		.PKT_TRANS_READ            (61),
		.PKT_TRANS_LOCK            (62),
		.PKT_SRC_ID_H              (85),
		.PKT_SRC_ID_L              (79),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (86),
		.PKT_BURSTWRAP_H           (69),
		.PKT_BURSTWRAP_L           (67),
		.PKT_BYTE_CNT_H            (66),
		.PKT_BYTE_CNT_L            (64),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (72),
		.PKT_BURST_SIZE_L          (70),
		.ST_CHANNEL_W              (99),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) ch0_yn1_l_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                           //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                //       clk_reset.reset
		.m0_address              (ch0_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ch0_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ch0_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ch0_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ch0_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ch0_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ch0_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ch0_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ch0_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ch0_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ch0_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ch0_yn1_l_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ch0_yn1_l_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ch0_yn1_l_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ch0_yn1_l_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ch0_yn1_l_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src18_ready),                                                    //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src18_valid),                                                    //                .valid
		.cp_data                 (cmd_xbar_demux_001_src18_data),                                                     //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src18_startofpacket),                                            //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src18_endofpacket),                                              //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src18_channel),                                                  //                .channel
		.rf_sink_ready           (ch0_yn1_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ch0_yn1_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ch0_yn1_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ch0_yn1_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ch0_yn1_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ch0_yn1_l_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ch0_yn1_l_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ch0_yn1_l_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ch0_yn1_l_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ch0_yn1_l_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ch0_yn1_l_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ch0_yn1_l_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (ch0_yn1_l_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (ch0_yn1_l_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ch0_yn1_l_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ch0_yn1_l_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                             //     (terminated)
		.m0_writeresponserequest (),                                                                                  //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                               //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ch0_yn1_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                           //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                // clk_reset.reset
		.in_data           (ch0_yn1_l_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ch0_yn1_l_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ch0_yn1_l_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ch0_yn1_l_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ch0_yn1_l_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ch0_yn1_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ch0_yn1_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ch0_yn1_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ch0_yn1_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ch0_yn1_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                             // (terminated)
		.csr_read          (1'b0),                                                                              // (terminated)
		.csr_write         (1'b0),                                                                              // (terminated)
		.csr_readdata      (),                                                                                  // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                              // (terminated)
		.almost_full_data  (),                                                                                  // (terminated)
		.almost_empty_data (),                                                                                  // (terminated)
		.in_empty          (1'b0),                                                                              // (terminated)
		.out_empty         (),                                                                                  // (terminated)
		.in_error          (1'b0),                                                                              // (terminated)
		.out_error         (),                                                                                  // (terminated)
		.in_channel        (1'b0),                                                                              // (terminated)
		.out_channel       ()                                                                                   // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (77),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (57),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (58),
		.PKT_TRANS_POSTED          (59),
		.PKT_TRANS_WRITE           (60),
		.PKT_TRANS_READ            (61),
		.PKT_TRANS_LOCK            (62),
		.PKT_SRC_ID_H              (85),
		.PKT_SRC_ID_L              (79),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (86),
		.PKT_BURSTWRAP_H           (69),
		.PKT_BURSTWRAP_L           (67),
		.PKT_BYTE_CNT_H            (66),
		.PKT_BYTE_CNT_L            (64),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (72),
		.PKT_BURST_SIZE_L          (70),
		.ST_CHANNEL_W              (99),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) ch0_yn1_ml_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                            //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                 //       clk_reset.reset
		.m0_address              (ch0_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ch0_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ch0_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ch0_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ch0_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ch0_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ch0_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ch0_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ch0_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ch0_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ch0_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ch0_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ch0_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ch0_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ch0_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ch0_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src19_ready),                                                     //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src19_valid),                                                     //                .valid
		.cp_data                 (cmd_xbar_demux_001_src19_data),                                                      //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src19_startofpacket),                                             //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src19_endofpacket),                                               //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src19_channel),                                                   //                .channel
		.rf_sink_ready           (ch0_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ch0_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ch0_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ch0_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ch0_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ch0_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ch0_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ch0_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ch0_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ch0_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ch0_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ch0_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (ch0_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (ch0_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ch0_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ch0_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                              //     (terminated)
		.m0_writeresponserequest (),                                                                                   //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ch0_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                            //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                 // clk_reset.reset
		.in_data           (ch0_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ch0_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ch0_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ch0_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ch0_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ch0_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ch0_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ch0_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ch0_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ch0_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                              // (terminated)
		.csr_read          (1'b0),                                                                               // (terminated)
		.csr_write         (1'b0),                                                                               // (terminated)
		.csr_readdata      (),                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                               // (terminated)
		.almost_full_data  (),                                                                                   // (terminated)
		.almost_empty_data (),                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                               // (terminated)
		.out_empty         (),                                                                                   // (terminated)
		.in_error          (1'b0),                                                                               // (terminated)
		.out_error         (),                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                               // (terminated)
		.out_channel       ()                                                                                    // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (77),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (57),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (58),
		.PKT_TRANS_POSTED          (59),
		.PKT_TRANS_WRITE           (60),
		.PKT_TRANS_READ            (61),
		.PKT_TRANS_LOCK            (62),
		.PKT_SRC_ID_H              (85),
		.PKT_SRC_ID_L              (79),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (86),
		.PKT_BURSTWRAP_H           (69),
		.PKT_BURSTWRAP_L           (67),
		.PKT_BYTE_CNT_H            (66),
		.PKT_BYTE_CNT_L            (64),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (72),
		.PKT_BURST_SIZE_L          (70),
		.ST_CHANNEL_W              (99),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) ch0_yn1_mu_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                            //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                 //       clk_reset.reset
		.m0_address              (ch0_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ch0_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ch0_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ch0_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ch0_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ch0_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ch0_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ch0_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ch0_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ch0_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ch0_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ch0_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ch0_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ch0_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ch0_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ch0_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src20_ready),                                                     //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src20_valid),                                                     //                .valid
		.cp_data                 (cmd_xbar_demux_001_src20_data),                                                      //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src20_startofpacket),                                             //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src20_endofpacket),                                               //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src20_channel),                                                   //                .channel
		.rf_sink_ready           (ch0_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ch0_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ch0_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ch0_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ch0_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ch0_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ch0_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ch0_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ch0_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ch0_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ch0_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ch0_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (ch0_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (ch0_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ch0_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ch0_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                              //     (terminated)
		.m0_writeresponserequest (),                                                                                   //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ch0_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                            //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                 // clk_reset.reset
		.in_data           (ch0_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ch0_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ch0_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ch0_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ch0_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ch0_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ch0_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ch0_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ch0_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ch0_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                              // (terminated)
		.csr_read          (1'b0),                                                                               // (terminated)
		.csr_write         (1'b0),                                                                               // (terminated)
		.csr_readdata      (),                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                               // (terminated)
		.almost_full_data  (),                                                                                   // (terminated)
		.almost_empty_data (),                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                               // (terminated)
		.out_empty         (),                                                                                   // (terminated)
		.in_error          (1'b0),                                                                               // (terminated)
		.out_error         (),                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                               // (terminated)
		.out_channel       ()                                                                                    // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (77),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (57),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (58),
		.PKT_TRANS_POSTED          (59),
		.PKT_TRANS_WRITE           (60),
		.PKT_TRANS_READ            (61),
		.PKT_TRANS_LOCK            (62),
		.PKT_SRC_ID_H              (85),
		.PKT_SRC_ID_L              (79),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (86),
		.PKT_BURSTWRAP_H           (69),
		.PKT_BURSTWRAP_L           (67),
		.PKT_BYTE_CNT_H            (66),
		.PKT_BYTE_CNT_L            (64),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (72),
		.PKT_BURST_SIZE_L          (70),
		.ST_CHANNEL_W              (99),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) ch0_yn1_u_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                           //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                //       clk_reset.reset
		.m0_address              (ch0_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ch0_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ch0_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ch0_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ch0_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ch0_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ch0_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ch0_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ch0_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ch0_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ch0_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ch0_yn1_u_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ch0_yn1_u_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ch0_yn1_u_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ch0_yn1_u_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ch0_yn1_u_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src21_ready),                                                    //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src21_valid),                                                    //                .valid
		.cp_data                 (cmd_xbar_demux_001_src21_data),                                                     //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src21_startofpacket),                                            //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src21_endofpacket),                                              //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src21_channel),                                                  //                .channel
		.rf_sink_ready           (ch0_yn1_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ch0_yn1_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ch0_yn1_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ch0_yn1_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ch0_yn1_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ch0_yn1_u_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ch0_yn1_u_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ch0_yn1_u_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ch0_yn1_u_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ch0_yn1_u_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ch0_yn1_u_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ch0_yn1_u_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (ch0_yn1_u_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (ch0_yn1_u_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ch0_yn1_u_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ch0_yn1_u_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                             //     (terminated)
		.m0_writeresponserequest (),                                                                                  //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                               //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ch0_yn1_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                           //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                // clk_reset.reset
		.in_data           (ch0_yn1_u_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ch0_yn1_u_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ch0_yn1_u_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ch0_yn1_u_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ch0_yn1_u_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ch0_yn1_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ch0_yn1_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ch0_yn1_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ch0_yn1_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ch0_yn1_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                             // (terminated)
		.csr_read          (1'b0),                                                                              // (terminated)
		.csr_write         (1'b0),                                                                              // (terminated)
		.csr_readdata      (),                                                                                  // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                              // (terminated)
		.almost_full_data  (),                                                                                  // (terminated)
		.almost_empty_data (),                                                                                  // (terminated)
		.in_empty          (1'b0),                                                                              // (terminated)
		.out_empty         (),                                                                                  // (terminated)
		.in_error          (1'b0),                                                                              // (terminated)
		.out_error         (),                                                                                  // (terminated)
		.in_channel        (1'b0),                                                                              // (terminated)
		.out_channel       ()                                                                                   // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (77),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (57),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (58),
		.PKT_TRANS_POSTED          (59),
		.PKT_TRANS_WRITE           (60),
		.PKT_TRANS_READ            (61),
		.PKT_TRANS_LOCK            (62),
		.PKT_SRC_ID_H              (85),
		.PKT_SRC_ID_L              (79),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (86),
		.PKT_BURSTWRAP_H           (69),
		.PKT_BURSTWRAP_L           (67),
		.PKT_BYTE_CNT_H            (66),
		.PKT_BYTE_CNT_L            (64),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (72),
		.PKT_BURST_SIZE_L          (70),
		.ST_CHANNEL_W              (99),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) ch0_time_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                          //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                               //       clk_reset.reset
		.m0_address              (ch0_time_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ch0_time_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ch0_time_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ch0_time_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ch0_time_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ch0_time_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ch0_time_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ch0_time_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ch0_time_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ch0_time_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ch0_time_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ch0_time_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ch0_time_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ch0_time_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ch0_time_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ch0_time_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src22_ready),                                                   //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src22_valid),                                                   //                .valid
		.cp_data                 (cmd_xbar_demux_001_src22_data),                                                    //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src22_startofpacket),                                           //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src22_endofpacket),                                             //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src22_channel),                                                 //                .channel
		.rf_sink_ready           (ch0_time_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ch0_time_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ch0_time_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ch0_time_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ch0_time_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ch0_time_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ch0_time_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ch0_time_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ch0_time_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ch0_time_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ch0_time_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ch0_time_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (ch0_time_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (ch0_time_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ch0_time_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ch0_time_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                            //     (terminated)
		.m0_writeresponserequest (),                                                                                 //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                              //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ch0_time_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                          //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                               // clk_reset.reset
		.in_data           (ch0_time_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ch0_time_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ch0_time_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ch0_time_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ch0_time_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ch0_time_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ch0_time_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ch0_time_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ch0_time_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ch0_time_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                            // (terminated)
		.csr_read          (1'b0),                                                                             // (terminated)
		.csr_write         (1'b0),                                                                             // (terminated)
		.csr_readdata      (),                                                                                 // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                             // (terminated)
		.almost_full_data  (),                                                                                 // (terminated)
		.almost_empty_data (),                                                                                 // (terminated)
		.in_empty          (1'b0),                                                                             // (terminated)
		.out_empty         (),                                                                                 // (terminated)
		.in_error          (1'b0),                                                                             // (terminated)
		.out_error         (),                                                                                 // (terminated)
		.in_channel        (1'b0),                                                                             // (terminated)
		.out_channel       ()                                                                                  // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (77),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (57),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (58),
		.PKT_TRANS_POSTED          (59),
		.PKT_TRANS_WRITE           (60),
		.PKT_TRANS_READ            (61),
		.PKT_TRANS_LOCK            (62),
		.PKT_SRC_ID_H              (85),
		.PKT_SRC_ID_L              (79),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (86),
		.PKT_BURSTWRAP_H           (69),
		.PKT_BURSTWRAP_L           (67),
		.PKT_BYTE_CNT_H            (66),
		.PKT_BYTE_CNT_L            (64),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (72),
		.PKT_BURST_SIZE_L          (70),
		.ST_CHANNEL_W              (99),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) ch0_yn2_mu_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                            //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                 //       clk_reset.reset
		.m0_address              (ch0_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ch0_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ch0_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ch0_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ch0_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ch0_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ch0_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ch0_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ch0_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ch0_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ch0_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ch0_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ch0_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ch0_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ch0_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ch0_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src23_ready),                                                     //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src23_valid),                                                     //                .valid
		.cp_data                 (cmd_xbar_demux_001_src23_data),                                                      //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src23_startofpacket),                                             //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src23_endofpacket),                                               //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src23_channel),                                                   //                .channel
		.rf_sink_ready           (ch0_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ch0_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ch0_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ch0_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ch0_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ch0_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ch0_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ch0_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ch0_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ch0_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ch0_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ch0_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (ch0_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (ch0_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ch0_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ch0_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                              //     (terminated)
		.m0_writeresponserequest (),                                                                                   //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ch0_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                            //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                 // clk_reset.reset
		.in_data           (ch0_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ch0_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ch0_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ch0_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ch0_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ch0_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ch0_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ch0_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ch0_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ch0_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                              // (terminated)
		.csr_read          (1'b0),                                                                               // (terminated)
		.csr_write         (1'b0),                                                                               // (terminated)
		.csr_readdata      (),                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                               // (terminated)
		.almost_full_data  (),                                                                                   // (terminated)
		.almost_empty_data (),                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                               // (terminated)
		.out_empty         (),                                                                                   // (terminated)
		.in_error          (1'b0),                                                                               // (terminated)
		.out_error         (),                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                               // (terminated)
		.out_channel       ()                                                                                    // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (77),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (57),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (58),
		.PKT_TRANS_POSTED          (59),
		.PKT_TRANS_WRITE           (60),
		.PKT_TRANS_READ            (61),
		.PKT_TRANS_LOCK            (62),
		.PKT_SRC_ID_H              (85),
		.PKT_SRC_ID_L              (79),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (86),
		.PKT_BURSTWRAP_H           (69),
		.PKT_BURSTWRAP_L           (67),
		.PKT_BYTE_CNT_H            (66),
		.PKT_BYTE_CNT_L            (64),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (72),
		.PKT_BURST_SIZE_L          (70),
		.ST_CHANNEL_W              (99),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) ch0_yn2_ml_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                            //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                 //       clk_reset.reset
		.m0_address              (ch0_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ch0_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ch0_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ch0_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ch0_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ch0_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ch0_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ch0_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ch0_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ch0_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ch0_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ch0_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ch0_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ch0_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ch0_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ch0_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src24_ready),                                                     //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src24_valid),                                                     //                .valid
		.cp_data                 (cmd_xbar_demux_001_src24_data),                                                      //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src24_startofpacket),                                             //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src24_endofpacket),                                               //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src24_channel),                                                   //                .channel
		.rf_sink_ready           (ch0_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ch0_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ch0_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ch0_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ch0_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ch0_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ch0_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ch0_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ch0_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ch0_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ch0_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ch0_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (ch0_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (ch0_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ch0_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ch0_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                              //     (terminated)
		.m0_writeresponserequest (),                                                                                   //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ch0_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                            //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                 // clk_reset.reset
		.in_data           (ch0_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ch0_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ch0_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ch0_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ch0_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ch0_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ch0_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ch0_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ch0_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ch0_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                              // (terminated)
		.csr_read          (1'b0),                                                                               // (terminated)
		.csr_write         (1'b0),                                                                               // (terminated)
		.csr_readdata      (),                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                               // (terminated)
		.almost_full_data  (),                                                                                   // (terminated)
		.almost_empty_data (),                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                               // (terminated)
		.out_empty         (),                                                                                   // (terminated)
		.in_error          (1'b0),                                                                               // (terminated)
		.out_error         (),                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                               // (terminated)
		.out_channel       ()                                                                                    // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (77),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (57),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (58),
		.PKT_TRANS_POSTED          (59),
		.PKT_TRANS_WRITE           (60),
		.PKT_TRANS_READ            (61),
		.PKT_TRANS_LOCK            (62),
		.PKT_SRC_ID_H              (85),
		.PKT_SRC_ID_L              (79),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (86),
		.PKT_BURSTWRAP_H           (69),
		.PKT_BURSTWRAP_L           (67),
		.PKT_BYTE_CNT_H            (66),
		.PKT_BYTE_CNT_L            (64),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (72),
		.PKT_BURST_SIZE_L          (70),
		.ST_CHANNEL_W              (99),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) ch0_yn2_u_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                           //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                //       clk_reset.reset
		.m0_address              (ch0_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ch0_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ch0_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ch0_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ch0_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ch0_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ch0_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ch0_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ch0_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ch0_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ch0_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ch0_yn2_u_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ch0_yn2_u_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ch0_yn2_u_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ch0_yn2_u_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ch0_yn2_u_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src25_ready),                                                    //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src25_valid),                                                    //                .valid
		.cp_data                 (cmd_xbar_demux_001_src25_data),                                                     //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src25_startofpacket),                                            //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src25_endofpacket),                                              //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src25_channel),                                                  //                .channel
		.rf_sink_ready           (ch0_yn2_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ch0_yn2_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ch0_yn2_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ch0_yn2_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ch0_yn2_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ch0_yn2_u_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ch0_yn2_u_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ch0_yn2_u_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ch0_yn2_u_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ch0_yn2_u_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ch0_yn2_u_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ch0_yn2_u_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (ch0_yn2_u_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (ch0_yn2_u_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ch0_yn2_u_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ch0_yn2_u_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                             //     (terminated)
		.m0_writeresponserequest (),                                                                                  //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                               //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ch0_yn2_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                           //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                // clk_reset.reset
		.in_data           (ch0_yn2_u_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ch0_yn2_u_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ch0_yn2_u_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ch0_yn2_u_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ch0_yn2_u_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ch0_yn2_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ch0_yn2_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ch0_yn2_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ch0_yn2_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ch0_yn2_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                             // (terminated)
		.csr_read          (1'b0),                                                                              // (terminated)
		.csr_write         (1'b0),                                                                              // (terminated)
		.csr_readdata      (),                                                                                  // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                              // (terminated)
		.almost_full_data  (),                                                                                  // (terminated)
		.almost_empty_data (),                                                                                  // (terminated)
		.in_empty          (1'b0),                                                                              // (terminated)
		.out_empty         (),                                                                                  // (terminated)
		.in_error          (1'b0),                                                                              // (terminated)
		.out_error         (),                                                                                  // (terminated)
		.in_channel        (1'b0),                                                                              // (terminated)
		.out_channel       ()                                                                                   // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (77),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (57),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (58),
		.PKT_TRANS_POSTED          (59),
		.PKT_TRANS_WRITE           (60),
		.PKT_TRANS_READ            (61),
		.PKT_TRANS_LOCK            (62),
		.PKT_SRC_ID_H              (85),
		.PKT_SRC_ID_L              (79),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (86),
		.PKT_BURSTWRAP_H           (69),
		.PKT_BURSTWRAP_L           (67),
		.PKT_BYTE_CNT_H            (66),
		.PKT_BYTE_CNT_L            (64),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (72),
		.PKT_BURST_SIZE_L          (70),
		.ST_CHANNEL_W              (99),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) ch0_yn2_l_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                           //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                //       clk_reset.reset
		.m0_address              (ch0_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ch0_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ch0_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ch0_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ch0_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ch0_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ch0_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ch0_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ch0_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ch0_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ch0_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ch0_yn2_l_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ch0_yn2_l_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ch0_yn2_l_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ch0_yn2_l_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ch0_yn2_l_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src26_ready),                                                    //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src26_valid),                                                    //                .valid
		.cp_data                 (cmd_xbar_demux_001_src26_data),                                                     //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src26_startofpacket),                                            //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src26_endofpacket),                                              //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src26_channel),                                                  //                .channel
		.rf_sink_ready           (ch0_yn2_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ch0_yn2_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ch0_yn2_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ch0_yn2_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ch0_yn2_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ch0_yn2_l_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ch0_yn2_l_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ch0_yn2_l_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ch0_yn2_l_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ch0_yn2_l_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ch0_yn2_l_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ch0_yn2_l_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (ch0_yn2_l_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (ch0_yn2_l_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ch0_yn2_l_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ch0_yn2_l_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                             //     (terminated)
		.m0_writeresponserequest (),                                                                                  //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                               //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ch0_yn2_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                           //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                // clk_reset.reset
		.in_data           (ch0_yn2_l_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ch0_yn2_l_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ch0_yn2_l_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ch0_yn2_l_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ch0_yn2_l_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ch0_yn2_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ch0_yn2_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ch0_yn2_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ch0_yn2_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ch0_yn2_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                             // (terminated)
		.csr_read          (1'b0),                                                                              // (terminated)
		.csr_write         (1'b0),                                                                              // (terminated)
		.csr_readdata      (),                                                                                  // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                              // (terminated)
		.almost_full_data  (),                                                                                  // (terminated)
		.almost_empty_data (),                                                                                  // (terminated)
		.in_empty          (1'b0),                                                                              // (terminated)
		.out_empty         (),                                                                                  // (terminated)
		.in_error          (1'b0),                                                                              // (terminated)
		.out_error         (),                                                                                  // (terminated)
		.in_channel        (1'b0),                                                                              // (terminated)
		.out_channel       ()                                                                                   // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (77),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (57),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (58),
		.PKT_TRANS_POSTED          (59),
		.PKT_TRANS_WRITE           (60),
		.PKT_TRANS_READ            (61),
		.PKT_TRANS_LOCK            (62),
		.PKT_SRC_ID_H              (85),
		.PKT_SRC_ID_L              (79),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (86),
		.PKT_BURSTWRAP_H           (69),
		.PKT_BURSTWRAP_L           (67),
		.PKT_BYTE_CNT_H            (66),
		.PKT_BYTE_CNT_L            (64),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (72),
		.PKT_BURST_SIZE_L          (70),
		.ST_CHANNEL_W              (99),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) ch0_yn3_l_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                           //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                //       clk_reset.reset
		.m0_address              (ch0_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ch0_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ch0_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ch0_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ch0_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ch0_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ch0_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ch0_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ch0_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ch0_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ch0_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ch0_yn3_l_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ch0_yn3_l_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ch0_yn3_l_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ch0_yn3_l_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ch0_yn3_l_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src27_ready),                                                    //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src27_valid),                                                    //                .valid
		.cp_data                 (cmd_xbar_demux_001_src27_data),                                                     //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src27_startofpacket),                                            //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src27_endofpacket),                                              //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src27_channel),                                                  //                .channel
		.rf_sink_ready           (ch0_yn3_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ch0_yn3_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ch0_yn3_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ch0_yn3_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ch0_yn3_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ch0_yn3_l_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ch0_yn3_l_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ch0_yn3_l_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ch0_yn3_l_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ch0_yn3_l_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ch0_yn3_l_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ch0_yn3_l_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (ch0_yn3_l_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (ch0_yn3_l_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ch0_yn3_l_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ch0_yn3_l_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                             //     (terminated)
		.m0_writeresponserequest (),                                                                                  //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                               //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ch0_yn3_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                           //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                // clk_reset.reset
		.in_data           (ch0_yn3_l_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ch0_yn3_l_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ch0_yn3_l_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ch0_yn3_l_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ch0_yn3_l_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ch0_yn3_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ch0_yn3_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ch0_yn3_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ch0_yn3_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ch0_yn3_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                             // (terminated)
		.csr_read          (1'b0),                                                                              // (terminated)
		.csr_write         (1'b0),                                                                              // (terminated)
		.csr_readdata      (),                                                                                  // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                              // (terminated)
		.almost_full_data  (),                                                                                  // (terminated)
		.almost_empty_data (),                                                                                  // (terminated)
		.in_empty          (1'b0),                                                                              // (terminated)
		.out_empty         (),                                                                                  // (terminated)
		.in_error          (1'b0),                                                                              // (terminated)
		.out_error         (),                                                                                  // (terminated)
		.in_channel        (1'b0),                                                                              // (terminated)
		.out_channel       ()                                                                                   // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (77),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (57),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (58),
		.PKT_TRANS_POSTED          (59),
		.PKT_TRANS_WRITE           (60),
		.PKT_TRANS_READ            (61),
		.PKT_TRANS_LOCK            (62),
		.PKT_SRC_ID_H              (85),
		.PKT_SRC_ID_L              (79),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (86),
		.PKT_BURSTWRAP_H           (69),
		.PKT_BURSTWRAP_L           (67),
		.PKT_BYTE_CNT_H            (66),
		.PKT_BYTE_CNT_L            (64),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (72),
		.PKT_BURST_SIZE_L          (70),
		.ST_CHANNEL_W              (99),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) ch0_yn3_ml_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                            //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                 //       clk_reset.reset
		.m0_address              (ch0_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ch0_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ch0_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ch0_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ch0_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ch0_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ch0_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ch0_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ch0_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ch0_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ch0_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ch0_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ch0_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ch0_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ch0_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ch0_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src28_ready),                                                     //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src28_valid),                                                     //                .valid
		.cp_data                 (cmd_xbar_demux_001_src28_data),                                                      //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src28_startofpacket),                                             //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src28_endofpacket),                                               //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src28_channel),                                                   //                .channel
		.rf_sink_ready           (ch0_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ch0_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ch0_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ch0_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ch0_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ch0_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ch0_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ch0_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ch0_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ch0_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ch0_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ch0_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (ch0_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (ch0_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ch0_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ch0_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                              //     (terminated)
		.m0_writeresponserequest (),                                                                                   //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ch0_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                            //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                 // clk_reset.reset
		.in_data           (ch0_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ch0_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ch0_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ch0_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ch0_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ch0_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ch0_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ch0_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ch0_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ch0_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                              // (terminated)
		.csr_read          (1'b0),                                                                               // (terminated)
		.csr_write         (1'b0),                                                                               // (terminated)
		.csr_readdata      (),                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                               // (terminated)
		.almost_full_data  (),                                                                                   // (terminated)
		.almost_empty_data (),                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                               // (terminated)
		.out_empty         (),                                                                                   // (terminated)
		.in_error          (1'b0),                                                                               // (terminated)
		.out_error         (),                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                               // (terminated)
		.out_channel       ()                                                                                    // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (77),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (57),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (58),
		.PKT_TRANS_POSTED          (59),
		.PKT_TRANS_WRITE           (60),
		.PKT_TRANS_READ            (61),
		.PKT_TRANS_LOCK            (62),
		.PKT_SRC_ID_H              (85),
		.PKT_SRC_ID_L              (79),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (86),
		.PKT_BURSTWRAP_H           (69),
		.PKT_BURSTWRAP_L           (67),
		.PKT_BYTE_CNT_H            (66),
		.PKT_BYTE_CNT_L            (64),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (72),
		.PKT_BURST_SIZE_L          (70),
		.ST_CHANNEL_W              (99),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) ch0_yn3_mu_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                            //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                 //       clk_reset.reset
		.m0_address              (ch0_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ch0_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ch0_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ch0_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ch0_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ch0_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ch0_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ch0_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ch0_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ch0_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ch0_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ch0_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ch0_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ch0_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ch0_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ch0_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src29_ready),                                                     //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src29_valid),                                                     //                .valid
		.cp_data                 (cmd_xbar_demux_001_src29_data),                                                      //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src29_startofpacket),                                             //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src29_endofpacket),                                               //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src29_channel),                                                   //                .channel
		.rf_sink_ready           (ch0_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ch0_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ch0_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ch0_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ch0_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ch0_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ch0_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ch0_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ch0_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ch0_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ch0_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ch0_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (ch0_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (ch0_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ch0_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ch0_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                              //     (terminated)
		.m0_writeresponserequest (),                                                                                   //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ch0_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                            //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                 // clk_reset.reset
		.in_data           (ch0_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ch0_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ch0_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ch0_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ch0_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ch0_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ch0_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ch0_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ch0_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ch0_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                              // (terminated)
		.csr_read          (1'b0),                                                                               // (terminated)
		.csr_write         (1'b0),                                                                               // (terminated)
		.csr_readdata      (),                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                               // (terminated)
		.almost_full_data  (),                                                                                   // (terminated)
		.almost_empty_data (),                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                               // (terminated)
		.out_empty         (),                                                                                   // (terminated)
		.in_error          (1'b0),                                                                               // (terminated)
		.out_error         (),                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                               // (terminated)
		.out_channel       ()                                                                                    // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (77),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (57),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (58),
		.PKT_TRANS_POSTED          (59),
		.PKT_TRANS_WRITE           (60),
		.PKT_TRANS_READ            (61),
		.PKT_TRANS_LOCK            (62),
		.PKT_SRC_ID_H              (85),
		.PKT_SRC_ID_L              (79),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (86),
		.PKT_BURSTWRAP_H           (69),
		.PKT_BURSTWRAP_L           (67),
		.PKT_BYTE_CNT_H            (66),
		.PKT_BYTE_CNT_L            (64),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (72),
		.PKT_BURST_SIZE_L          (70),
		.ST_CHANNEL_W              (99),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) ch0_yn3_u_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                           //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                //       clk_reset.reset
		.m0_address              (ch0_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ch0_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ch0_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ch0_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ch0_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ch0_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ch0_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ch0_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ch0_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ch0_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ch0_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ch0_yn3_u_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ch0_yn3_u_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ch0_yn3_u_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ch0_yn3_u_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ch0_yn3_u_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src30_ready),                                                    //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src30_valid),                                                    //                .valid
		.cp_data                 (cmd_xbar_demux_001_src30_data),                                                     //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src30_startofpacket),                                            //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src30_endofpacket),                                              //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src30_channel),                                                  //                .channel
		.rf_sink_ready           (ch0_yn3_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ch0_yn3_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ch0_yn3_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ch0_yn3_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ch0_yn3_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ch0_yn3_u_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ch0_yn3_u_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ch0_yn3_u_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ch0_yn3_u_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ch0_yn3_u_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ch0_yn3_u_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ch0_yn3_u_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (ch0_yn3_u_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (ch0_yn3_u_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ch0_yn3_u_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ch0_yn3_u_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                             //     (terminated)
		.m0_writeresponserequest (),                                                                                  //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                               //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ch0_yn3_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                           //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                // clk_reset.reset
		.in_data           (ch0_yn3_u_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ch0_yn3_u_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ch0_yn3_u_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ch0_yn3_u_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ch0_yn3_u_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ch0_yn3_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ch0_yn3_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ch0_yn3_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ch0_yn3_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ch0_yn3_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                             // (terminated)
		.csr_read          (1'b0),                                                                              // (terminated)
		.csr_write         (1'b0),                                                                              // (terminated)
		.csr_readdata      (),                                                                                  // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                              // (terminated)
		.almost_full_data  (),                                                                                  // (terminated)
		.almost_empty_data (),                                                                                  // (terminated)
		.in_empty          (1'b0),                                                                              // (terminated)
		.out_empty         (),                                                                                  // (terminated)
		.in_error          (1'b0),                                                                              // (terminated)
		.out_error         (),                                                                                  // (terminated)
		.in_channel        (1'b0),                                                                              // (terminated)
		.out_channel       ()                                                                                   // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (77),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (57),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (58),
		.PKT_TRANS_POSTED          (59),
		.PKT_TRANS_WRITE           (60),
		.PKT_TRANS_READ            (61),
		.PKT_TRANS_LOCK            (62),
		.PKT_SRC_ID_H              (85),
		.PKT_SRC_ID_L              (79),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (86),
		.PKT_BURSTWRAP_H           (69),
		.PKT_BURSTWRAP_L           (67),
		.PKT_BYTE_CNT_H            (66),
		.PKT_BYTE_CNT_L            (64),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (72),
		.PKT_BURST_SIZE_L          (70),
		.ST_CHANNEL_W              (99),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) ch1_timer_rst_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                               //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                    //       clk_reset.reset
		.m0_address              (ch1_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ch1_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ch1_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ch1_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ch1_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ch1_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ch1_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ch1_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ch1_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ch1_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ch1_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ch1_timer_rst_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ch1_timer_rst_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ch1_timer_rst_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ch1_timer_rst_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ch1_timer_rst_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src31_ready),                                                        //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src31_valid),                                                        //                .valid
		.cp_data                 (cmd_xbar_demux_001_src31_data),                                                         //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src31_startofpacket),                                                //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src31_endofpacket),                                                  //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src31_channel),                                                      //                .channel
		.rf_sink_ready           (ch1_timer_rst_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ch1_timer_rst_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ch1_timer_rst_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ch1_timer_rst_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ch1_timer_rst_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ch1_timer_rst_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ch1_timer_rst_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ch1_timer_rst_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ch1_timer_rst_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ch1_timer_rst_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ch1_timer_rst_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ch1_timer_rst_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (ch1_timer_rst_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (ch1_timer_rst_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ch1_timer_rst_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ch1_timer_rst_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                 //     (terminated)
		.m0_writeresponserequest (),                                                                                      //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                   //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ch1_timer_rst_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                               //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                    // clk_reset.reset
		.in_data           (ch1_timer_rst_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ch1_timer_rst_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ch1_timer_rst_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ch1_timer_rst_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ch1_timer_rst_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ch1_timer_rst_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ch1_timer_rst_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ch1_timer_rst_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ch1_timer_rst_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ch1_timer_rst_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                 // (terminated)
		.csr_read          (1'b0),                                                                                  // (terminated)
		.csr_write         (1'b0),                                                                                  // (terminated)
		.csr_readdata      (),                                                                                      // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                  // (terminated)
		.almost_full_data  (),                                                                                      // (terminated)
		.almost_empty_data (),                                                                                      // (terminated)
		.in_empty          (1'b0),                                                                                  // (terminated)
		.out_empty         (),                                                                                      // (terminated)
		.in_error          (1'b0),                                                                                  // (terminated)
		.out_error         (),                                                                                      // (terminated)
		.in_channel        (1'b0),                                                                                  // (terminated)
		.out_channel       ()                                                                                       // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (77),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (57),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (58),
		.PKT_TRANS_POSTED          (59),
		.PKT_TRANS_WRITE           (60),
		.PKT_TRANS_READ            (61),
		.PKT_TRANS_LOCK            (62),
		.PKT_SRC_ID_H              (85),
		.PKT_SRC_ID_L              (79),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (86),
		.PKT_BURSTWRAP_H           (69),
		.PKT_BURSTWRAP_L           (67),
		.PKT_BYTE_CNT_H            (66),
		.PKT_BYTE_CNT_L            (64),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (72),
		.PKT_BURST_SIZE_L          (70),
		.ST_CHANNEL_W              (99),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) ch1_thresh_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                            //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                 //       clk_reset.reset
		.m0_address              (ch1_thresh_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ch1_thresh_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ch1_thresh_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ch1_thresh_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ch1_thresh_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ch1_thresh_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ch1_thresh_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ch1_thresh_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ch1_thresh_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ch1_thresh_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ch1_thresh_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ch1_thresh_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ch1_thresh_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ch1_thresh_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ch1_thresh_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ch1_thresh_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src32_ready),                                                     //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src32_valid),                                                     //                .valid
		.cp_data                 (cmd_xbar_demux_001_src32_data),                                                      //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src32_startofpacket),                                             //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src32_endofpacket),                                               //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src32_channel),                                                   //                .channel
		.rf_sink_ready           (ch1_thresh_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ch1_thresh_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ch1_thresh_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ch1_thresh_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ch1_thresh_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ch1_thresh_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ch1_thresh_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ch1_thresh_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ch1_thresh_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ch1_thresh_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ch1_thresh_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ch1_thresh_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (ch1_thresh_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (ch1_thresh_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ch1_thresh_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ch1_thresh_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                              //     (terminated)
		.m0_writeresponserequest (),                                                                                   //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ch1_thresh_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                            //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                 // clk_reset.reset
		.in_data           (ch1_thresh_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ch1_thresh_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ch1_thresh_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ch1_thresh_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ch1_thresh_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ch1_thresh_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ch1_thresh_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ch1_thresh_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ch1_thresh_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ch1_thresh_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                              // (terminated)
		.csr_read          (1'b0),                                                                               // (terminated)
		.csr_write         (1'b0),                                                                               // (terminated)
		.csr_readdata      (),                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                               // (terminated)
		.almost_full_data  (),                                                                                   // (terminated)
		.almost_empty_data (),                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                               // (terminated)
		.out_empty         (),                                                                                   // (terminated)
		.in_error          (1'b0),                                                                               // (terminated)
		.out_error         (),                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                               // (terminated)
		.out_channel       ()                                                                                    // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (77),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (57),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (58),
		.PKT_TRANS_POSTED          (59),
		.PKT_TRANS_WRITE           (60),
		.PKT_TRANS_READ            (61),
		.PKT_TRANS_LOCK            (62),
		.PKT_SRC_ID_H              (85),
		.PKT_SRC_ID_L              (79),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (86),
		.PKT_BURSTWRAP_H           (69),
		.PKT_BURSTWRAP_L           (67),
		.PKT_BYTE_CNT_H            (66),
		.PKT_BYTE_CNT_L            (64),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (72),
		.PKT_BURST_SIZE_L          (70),
		.ST_CHANNEL_W              (99),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) ch1_rd_peak_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                             //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                  //       clk_reset.reset
		.m0_address              (ch1_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ch1_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ch1_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ch1_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ch1_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ch1_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ch1_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ch1_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ch1_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ch1_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ch1_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ch1_rd_peak_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ch1_rd_peak_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ch1_rd_peak_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ch1_rd_peak_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ch1_rd_peak_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src33_ready),                                                      //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src33_valid),                                                      //                .valid
		.cp_data                 (cmd_xbar_demux_001_src33_data),                                                       //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src33_startofpacket),                                              //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src33_endofpacket),                                                //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src33_channel),                                                    //                .channel
		.rf_sink_ready           (ch1_rd_peak_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ch1_rd_peak_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ch1_rd_peak_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ch1_rd_peak_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ch1_rd_peak_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ch1_rd_peak_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ch1_rd_peak_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ch1_rd_peak_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ch1_rd_peak_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ch1_rd_peak_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ch1_rd_peak_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ch1_rd_peak_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (ch1_rd_peak_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (ch1_rd_peak_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ch1_rd_peak_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ch1_rd_peak_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                               //     (terminated)
		.m0_writeresponserequest (),                                                                                    //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                 //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ch1_rd_peak_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                             //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                  // clk_reset.reset
		.in_data           (ch1_rd_peak_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ch1_rd_peak_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ch1_rd_peak_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ch1_rd_peak_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ch1_rd_peak_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ch1_rd_peak_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ch1_rd_peak_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ch1_rd_peak_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ch1_rd_peak_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ch1_rd_peak_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                               // (terminated)
		.csr_read          (1'b0),                                                                                // (terminated)
		.csr_write         (1'b0),                                                                                // (terminated)
		.csr_readdata      (),                                                                                    // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                // (terminated)
		.almost_full_data  (),                                                                                    // (terminated)
		.almost_empty_data (),                                                                                    // (terminated)
		.in_empty          (1'b0),                                                                                // (terminated)
		.out_empty         (),                                                                                    // (terminated)
		.in_error          (1'b0),                                                                                // (terminated)
		.out_error         (),                                                                                    // (terminated)
		.in_channel        (1'b0),                                                                                // (terminated)
		.out_channel       ()                                                                                     // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (77),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (57),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (58),
		.PKT_TRANS_POSTED          (59),
		.PKT_TRANS_WRITE           (60),
		.PKT_TRANS_READ            (61),
		.PKT_TRANS_LOCK            (62),
		.PKT_SRC_ID_H              (85),
		.PKT_SRC_ID_L              (79),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (86),
		.PKT_BURSTWRAP_H           (69),
		.PKT_BURSTWRAP_L           (67),
		.PKT_BYTE_CNT_H            (66),
		.PKT_BYTE_CNT_L            (64),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (72),
		.PKT_BURST_SIZE_L          (70),
		.ST_CHANNEL_W              (99),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) ch1_peak_found_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                     //       clk_reset.reset
		.m0_address              (ch1_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ch1_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ch1_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ch1_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ch1_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ch1_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ch1_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ch1_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ch1_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ch1_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ch1_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ch1_peak_found_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ch1_peak_found_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ch1_peak_found_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ch1_peak_found_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ch1_peak_found_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src34_ready),                                                         //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src34_valid),                                                         //                .valid
		.cp_data                 (cmd_xbar_demux_001_src34_data),                                                          //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src34_startofpacket),                                                 //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src34_endofpacket),                                                   //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src34_channel),                                                       //                .channel
		.rf_sink_ready           (ch1_peak_found_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ch1_peak_found_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ch1_peak_found_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ch1_peak_found_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ch1_peak_found_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ch1_peak_found_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ch1_peak_found_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ch1_peak_found_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ch1_peak_found_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ch1_peak_found_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ch1_peak_found_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ch1_peak_found_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (ch1_peak_found_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (ch1_peak_found_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ch1_peak_found_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ch1_peak_found_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                  //     (terminated)
		.m0_writeresponserequest (),                                                                                       //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                    //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ch1_peak_found_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                     // clk_reset.reset
		.in_data           (ch1_peak_found_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ch1_peak_found_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ch1_peak_found_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ch1_peak_found_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ch1_peak_found_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ch1_peak_found_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ch1_peak_found_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ch1_peak_found_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ch1_peak_found_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ch1_peak_found_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                  // (terminated)
		.csr_read          (1'b0),                                                                                   // (terminated)
		.csr_write         (1'b0),                                                                                   // (terminated)
		.csr_readdata      (),                                                                                       // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                   // (terminated)
		.almost_full_data  (),                                                                                       // (terminated)
		.almost_empty_data (),                                                                                       // (terminated)
		.in_empty          (1'b0),                                                                                   // (terminated)
		.out_empty         (),                                                                                       // (terminated)
		.in_error          (1'b0),                                                                                   // (terminated)
		.out_error         (),                                                                                       // (terminated)
		.in_channel        (1'b0),                                                                                   // (terminated)
		.out_channel       ()                                                                                        // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (77),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (57),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (58),
		.PKT_TRANS_POSTED          (59),
		.PKT_TRANS_WRITE           (60),
		.PKT_TRANS_READ            (61),
		.PKT_TRANS_LOCK            (62),
		.PKT_SRC_ID_H              (85),
		.PKT_SRC_ID_L              (79),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (86),
		.PKT_BURSTWRAP_H           (69),
		.PKT_BURSTWRAP_L           (67),
		.PKT_BYTE_CNT_H            (66),
		.PKT_BYTE_CNT_L            (64),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (72),
		.PKT_BURST_SIZE_L          (70),
		.ST_CHANNEL_W              (99),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) ch1_time_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                          //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                               //       clk_reset.reset
		.m0_address              (ch1_time_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ch1_time_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ch1_time_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ch1_time_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ch1_time_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ch1_time_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ch1_time_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ch1_time_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ch1_time_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ch1_time_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ch1_time_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ch1_time_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ch1_time_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ch1_time_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ch1_time_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ch1_time_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src35_ready),                                                   //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src35_valid),                                                   //                .valid
		.cp_data                 (cmd_xbar_demux_001_src35_data),                                                    //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src35_startofpacket),                                           //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src35_endofpacket),                                             //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src35_channel),                                                 //                .channel
		.rf_sink_ready           (ch1_time_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ch1_time_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ch1_time_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ch1_time_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ch1_time_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ch1_time_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ch1_time_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ch1_time_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ch1_time_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ch1_time_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ch1_time_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ch1_time_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (ch1_time_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (ch1_time_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ch1_time_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ch1_time_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                            //     (terminated)
		.m0_writeresponserequest (),                                                                                 //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                              //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ch1_time_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                          //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                               // clk_reset.reset
		.in_data           (ch1_time_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ch1_time_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ch1_time_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ch1_time_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ch1_time_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ch1_time_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ch1_time_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ch1_time_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ch1_time_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ch1_time_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                            // (terminated)
		.csr_read          (1'b0),                                                                             // (terminated)
		.csr_write         (1'b0),                                                                             // (terminated)
		.csr_readdata      (),                                                                                 // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                             // (terminated)
		.almost_full_data  (),                                                                                 // (terminated)
		.almost_empty_data (),                                                                                 // (terminated)
		.in_empty          (1'b0),                                                                             // (terminated)
		.out_empty         (),                                                                                 // (terminated)
		.in_error          (1'b0),                                                                             // (terminated)
		.out_error         (),                                                                                 // (terminated)
		.in_channel        (1'b0),                                                                             // (terminated)
		.out_channel       ()                                                                                  // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (77),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (57),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (58),
		.PKT_TRANS_POSTED          (59),
		.PKT_TRANS_WRITE           (60),
		.PKT_TRANS_READ            (61),
		.PKT_TRANS_LOCK            (62),
		.PKT_SRC_ID_H              (85),
		.PKT_SRC_ID_L              (79),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (86),
		.PKT_BURSTWRAP_H           (69),
		.PKT_BURSTWRAP_L           (67),
		.PKT_BYTE_CNT_H            (66),
		.PKT_BYTE_CNT_L            (64),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (72),
		.PKT_BURST_SIZE_L          (70),
		.ST_CHANNEL_W              (99),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) ch1_yn1_u_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                           //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                //       clk_reset.reset
		.m0_address              (ch1_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ch1_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ch1_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ch1_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ch1_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ch1_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ch1_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ch1_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ch1_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ch1_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ch1_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ch1_yn1_u_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ch1_yn1_u_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ch1_yn1_u_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ch1_yn1_u_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ch1_yn1_u_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src36_ready),                                                    //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src36_valid),                                                    //                .valid
		.cp_data                 (cmd_xbar_demux_001_src36_data),                                                     //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src36_startofpacket),                                            //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src36_endofpacket),                                              //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src36_channel),                                                  //                .channel
		.rf_sink_ready           (ch1_yn1_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ch1_yn1_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ch1_yn1_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ch1_yn1_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ch1_yn1_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ch1_yn1_u_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ch1_yn1_u_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ch1_yn1_u_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ch1_yn1_u_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ch1_yn1_u_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ch1_yn1_u_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ch1_yn1_u_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (ch1_yn1_u_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (ch1_yn1_u_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ch1_yn1_u_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ch1_yn1_u_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                             //     (terminated)
		.m0_writeresponserequest (),                                                                                  //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                               //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ch1_yn1_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                           //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                // clk_reset.reset
		.in_data           (ch1_yn1_u_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ch1_yn1_u_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ch1_yn1_u_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ch1_yn1_u_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ch1_yn1_u_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ch1_yn1_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ch1_yn1_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ch1_yn1_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ch1_yn1_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ch1_yn1_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                             // (terminated)
		.csr_read          (1'b0),                                                                              // (terminated)
		.csr_write         (1'b0),                                                                              // (terminated)
		.csr_readdata      (),                                                                                  // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                              // (terminated)
		.almost_full_data  (),                                                                                  // (terminated)
		.almost_empty_data (),                                                                                  // (terminated)
		.in_empty          (1'b0),                                                                              // (terminated)
		.out_empty         (),                                                                                  // (terminated)
		.in_error          (1'b0),                                                                              // (terminated)
		.out_error         (),                                                                                  // (terminated)
		.in_channel        (1'b0),                                                                              // (terminated)
		.out_channel       ()                                                                                   // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (77),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (57),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (58),
		.PKT_TRANS_POSTED          (59),
		.PKT_TRANS_WRITE           (60),
		.PKT_TRANS_READ            (61),
		.PKT_TRANS_LOCK            (62),
		.PKT_SRC_ID_H              (85),
		.PKT_SRC_ID_L              (79),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (86),
		.PKT_BURSTWRAP_H           (69),
		.PKT_BURSTWRAP_L           (67),
		.PKT_BYTE_CNT_H            (66),
		.PKT_BYTE_CNT_L            (64),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (72),
		.PKT_BURST_SIZE_L          (70),
		.ST_CHANNEL_W              (99),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) ch1_yn1_mu_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                            //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                 //       clk_reset.reset
		.m0_address              (ch1_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ch1_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ch1_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ch1_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ch1_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ch1_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ch1_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ch1_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ch1_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ch1_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ch1_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ch1_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ch1_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ch1_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ch1_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ch1_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src37_ready),                                                     //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src37_valid),                                                     //                .valid
		.cp_data                 (cmd_xbar_demux_001_src37_data),                                                      //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src37_startofpacket),                                             //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src37_endofpacket),                                               //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src37_channel),                                                   //                .channel
		.rf_sink_ready           (ch1_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ch1_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ch1_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ch1_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ch1_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ch1_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ch1_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ch1_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ch1_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ch1_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ch1_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ch1_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (ch1_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (ch1_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ch1_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ch1_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                              //     (terminated)
		.m0_writeresponserequest (),                                                                                   //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ch1_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                            //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                 // clk_reset.reset
		.in_data           (ch1_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ch1_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ch1_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ch1_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ch1_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ch1_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ch1_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ch1_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ch1_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ch1_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                              // (terminated)
		.csr_read          (1'b0),                                                                               // (terminated)
		.csr_write         (1'b0),                                                                               // (terminated)
		.csr_readdata      (),                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                               // (terminated)
		.almost_full_data  (),                                                                                   // (terminated)
		.almost_empty_data (),                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                               // (terminated)
		.out_empty         (),                                                                                   // (terminated)
		.in_error          (1'b0),                                                                               // (terminated)
		.out_error         (),                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                               // (terminated)
		.out_channel       ()                                                                                    // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (77),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (57),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (58),
		.PKT_TRANS_POSTED          (59),
		.PKT_TRANS_WRITE           (60),
		.PKT_TRANS_READ            (61),
		.PKT_TRANS_LOCK            (62),
		.PKT_SRC_ID_H              (85),
		.PKT_SRC_ID_L              (79),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (86),
		.PKT_BURSTWRAP_H           (69),
		.PKT_BURSTWRAP_L           (67),
		.PKT_BYTE_CNT_H            (66),
		.PKT_BYTE_CNT_L            (64),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (72),
		.PKT_BURST_SIZE_L          (70),
		.ST_CHANNEL_W              (99),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) ch1_yn1_ml_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                            //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                 //       clk_reset.reset
		.m0_address              (ch1_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ch1_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ch1_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ch1_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ch1_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ch1_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ch1_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ch1_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ch1_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ch1_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ch1_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ch1_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ch1_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ch1_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ch1_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ch1_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src38_ready),                                                     //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src38_valid),                                                     //                .valid
		.cp_data                 (cmd_xbar_demux_001_src38_data),                                                      //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src38_startofpacket),                                             //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src38_endofpacket),                                               //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src38_channel),                                                   //                .channel
		.rf_sink_ready           (ch1_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ch1_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ch1_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ch1_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ch1_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ch1_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ch1_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ch1_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ch1_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ch1_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ch1_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ch1_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (ch1_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (ch1_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ch1_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ch1_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                              //     (terminated)
		.m0_writeresponserequest (),                                                                                   //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ch1_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                            //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                 // clk_reset.reset
		.in_data           (ch1_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ch1_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ch1_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ch1_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ch1_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ch1_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ch1_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ch1_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ch1_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ch1_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                              // (terminated)
		.csr_read          (1'b0),                                                                               // (terminated)
		.csr_write         (1'b0),                                                                               // (terminated)
		.csr_readdata      (),                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                               // (terminated)
		.almost_full_data  (),                                                                                   // (terminated)
		.almost_empty_data (),                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                               // (terminated)
		.out_empty         (),                                                                                   // (terminated)
		.in_error          (1'b0),                                                                               // (terminated)
		.out_error         (),                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                               // (terminated)
		.out_channel       ()                                                                                    // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (77),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (57),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (58),
		.PKT_TRANS_POSTED          (59),
		.PKT_TRANS_WRITE           (60),
		.PKT_TRANS_READ            (61),
		.PKT_TRANS_LOCK            (62),
		.PKT_SRC_ID_H              (85),
		.PKT_SRC_ID_L              (79),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (86),
		.PKT_BURSTWRAP_H           (69),
		.PKT_BURSTWRAP_L           (67),
		.PKT_BYTE_CNT_H            (66),
		.PKT_BYTE_CNT_L            (64),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (72),
		.PKT_BURST_SIZE_L          (70),
		.ST_CHANNEL_W              (99),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) ch1_yn1_l_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                           //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                //       clk_reset.reset
		.m0_address              (ch1_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ch1_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ch1_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ch1_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ch1_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ch1_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ch1_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ch1_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ch1_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ch1_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ch1_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ch1_yn1_l_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ch1_yn1_l_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ch1_yn1_l_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ch1_yn1_l_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ch1_yn1_l_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src39_ready),                                                    //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src39_valid),                                                    //                .valid
		.cp_data                 (cmd_xbar_demux_001_src39_data),                                                     //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src39_startofpacket),                                            //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src39_endofpacket),                                              //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src39_channel),                                                  //                .channel
		.rf_sink_ready           (ch1_yn1_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ch1_yn1_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ch1_yn1_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ch1_yn1_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ch1_yn1_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ch1_yn1_l_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ch1_yn1_l_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ch1_yn1_l_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ch1_yn1_l_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ch1_yn1_l_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ch1_yn1_l_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ch1_yn1_l_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (ch1_yn1_l_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (ch1_yn1_l_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ch1_yn1_l_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ch1_yn1_l_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                             //     (terminated)
		.m0_writeresponserequest (),                                                                                  //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                               //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ch1_yn1_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                           //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                // clk_reset.reset
		.in_data           (ch1_yn1_l_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ch1_yn1_l_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ch1_yn1_l_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ch1_yn1_l_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ch1_yn1_l_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ch1_yn1_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ch1_yn1_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ch1_yn1_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ch1_yn1_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ch1_yn1_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                             // (terminated)
		.csr_read          (1'b0),                                                                              // (terminated)
		.csr_write         (1'b0),                                                                              // (terminated)
		.csr_readdata      (),                                                                                  // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                              // (terminated)
		.almost_full_data  (),                                                                                  // (terminated)
		.almost_empty_data (),                                                                                  // (terminated)
		.in_empty          (1'b0),                                                                              // (terminated)
		.out_empty         (),                                                                                  // (terminated)
		.in_error          (1'b0),                                                                              // (terminated)
		.out_error         (),                                                                                  // (terminated)
		.in_channel        (1'b0),                                                                              // (terminated)
		.out_channel       ()                                                                                   // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (77),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (57),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (58),
		.PKT_TRANS_POSTED          (59),
		.PKT_TRANS_WRITE           (60),
		.PKT_TRANS_READ            (61),
		.PKT_TRANS_LOCK            (62),
		.PKT_SRC_ID_H              (85),
		.PKT_SRC_ID_L              (79),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (86),
		.PKT_BURSTWRAP_H           (69),
		.PKT_BURSTWRAP_L           (67),
		.PKT_BYTE_CNT_H            (66),
		.PKT_BYTE_CNT_L            (64),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (72),
		.PKT_BURST_SIZE_L          (70),
		.ST_CHANNEL_W              (99),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) ch1_yn2_u_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                           //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                //       clk_reset.reset
		.m0_address              (ch1_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ch1_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ch1_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ch1_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ch1_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ch1_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ch1_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ch1_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ch1_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ch1_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ch1_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ch1_yn2_u_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ch1_yn2_u_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ch1_yn2_u_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ch1_yn2_u_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ch1_yn2_u_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src40_ready),                                                    //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src40_valid),                                                    //                .valid
		.cp_data                 (cmd_xbar_demux_001_src40_data),                                                     //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src40_startofpacket),                                            //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src40_endofpacket),                                              //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src40_channel),                                                  //                .channel
		.rf_sink_ready           (ch1_yn2_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ch1_yn2_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ch1_yn2_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ch1_yn2_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ch1_yn2_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ch1_yn2_u_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ch1_yn2_u_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ch1_yn2_u_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ch1_yn2_u_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ch1_yn2_u_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ch1_yn2_u_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ch1_yn2_u_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (ch1_yn2_u_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (ch1_yn2_u_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ch1_yn2_u_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ch1_yn2_u_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                             //     (terminated)
		.m0_writeresponserequest (),                                                                                  //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                               //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ch1_yn2_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                           //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                // clk_reset.reset
		.in_data           (ch1_yn2_u_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ch1_yn2_u_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ch1_yn2_u_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ch1_yn2_u_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ch1_yn2_u_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ch1_yn2_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ch1_yn2_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ch1_yn2_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ch1_yn2_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ch1_yn2_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                             // (terminated)
		.csr_read          (1'b0),                                                                              // (terminated)
		.csr_write         (1'b0),                                                                              // (terminated)
		.csr_readdata      (),                                                                                  // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                              // (terminated)
		.almost_full_data  (),                                                                                  // (terminated)
		.almost_empty_data (),                                                                                  // (terminated)
		.in_empty          (1'b0),                                                                              // (terminated)
		.out_empty         (),                                                                                  // (terminated)
		.in_error          (1'b0),                                                                              // (terminated)
		.out_error         (),                                                                                  // (terminated)
		.in_channel        (1'b0),                                                                              // (terminated)
		.out_channel       ()                                                                                   // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (77),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (57),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (58),
		.PKT_TRANS_POSTED          (59),
		.PKT_TRANS_WRITE           (60),
		.PKT_TRANS_READ            (61),
		.PKT_TRANS_LOCK            (62),
		.PKT_SRC_ID_H              (85),
		.PKT_SRC_ID_L              (79),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (86),
		.PKT_BURSTWRAP_H           (69),
		.PKT_BURSTWRAP_L           (67),
		.PKT_BYTE_CNT_H            (66),
		.PKT_BYTE_CNT_L            (64),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (72),
		.PKT_BURST_SIZE_L          (70),
		.ST_CHANNEL_W              (99),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) ch1_yn2_mu_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                            //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                 //       clk_reset.reset
		.m0_address              (ch1_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ch1_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ch1_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ch1_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ch1_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ch1_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ch1_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ch1_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ch1_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ch1_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ch1_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ch1_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ch1_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ch1_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ch1_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ch1_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src41_ready),                                                     //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src41_valid),                                                     //                .valid
		.cp_data                 (cmd_xbar_demux_001_src41_data),                                                      //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src41_startofpacket),                                             //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src41_endofpacket),                                               //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src41_channel),                                                   //                .channel
		.rf_sink_ready           (ch1_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ch1_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ch1_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ch1_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ch1_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ch1_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ch1_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ch1_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ch1_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ch1_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ch1_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ch1_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (ch1_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (ch1_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ch1_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ch1_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                              //     (terminated)
		.m0_writeresponserequest (),                                                                                   //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ch1_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                            //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                 // clk_reset.reset
		.in_data           (ch1_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ch1_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ch1_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ch1_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ch1_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ch1_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ch1_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ch1_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ch1_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ch1_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                              // (terminated)
		.csr_read          (1'b0),                                                                               // (terminated)
		.csr_write         (1'b0),                                                                               // (terminated)
		.csr_readdata      (),                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                               // (terminated)
		.almost_full_data  (),                                                                                   // (terminated)
		.almost_empty_data (),                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                               // (terminated)
		.out_empty         (),                                                                                   // (terminated)
		.in_error          (1'b0),                                                                               // (terminated)
		.out_error         (),                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                               // (terminated)
		.out_channel       ()                                                                                    // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (77),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (57),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (58),
		.PKT_TRANS_POSTED          (59),
		.PKT_TRANS_WRITE           (60),
		.PKT_TRANS_READ            (61),
		.PKT_TRANS_LOCK            (62),
		.PKT_SRC_ID_H              (85),
		.PKT_SRC_ID_L              (79),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (86),
		.PKT_BURSTWRAP_H           (69),
		.PKT_BURSTWRAP_L           (67),
		.PKT_BYTE_CNT_H            (66),
		.PKT_BYTE_CNT_L            (64),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (72),
		.PKT_BURST_SIZE_L          (70),
		.ST_CHANNEL_W              (99),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) ch1_yn2_ml_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                            //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                 //       clk_reset.reset
		.m0_address              (ch1_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ch1_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ch1_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ch1_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ch1_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ch1_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ch1_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ch1_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ch1_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ch1_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ch1_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ch1_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ch1_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ch1_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ch1_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ch1_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src42_ready),                                                     //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src42_valid),                                                     //                .valid
		.cp_data                 (cmd_xbar_demux_001_src42_data),                                                      //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src42_startofpacket),                                             //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src42_endofpacket),                                               //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src42_channel),                                                   //                .channel
		.rf_sink_ready           (ch1_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ch1_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ch1_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ch1_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ch1_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ch1_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ch1_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ch1_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ch1_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ch1_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ch1_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ch1_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (ch1_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (ch1_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ch1_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ch1_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                              //     (terminated)
		.m0_writeresponserequest (),                                                                                   //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ch1_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                            //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                 // clk_reset.reset
		.in_data           (ch1_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ch1_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ch1_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ch1_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ch1_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ch1_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ch1_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ch1_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ch1_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ch1_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                              // (terminated)
		.csr_read          (1'b0),                                                                               // (terminated)
		.csr_write         (1'b0),                                                                               // (terminated)
		.csr_readdata      (),                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                               // (terminated)
		.almost_full_data  (),                                                                                   // (terminated)
		.almost_empty_data (),                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                               // (terminated)
		.out_empty         (),                                                                                   // (terminated)
		.in_error          (1'b0),                                                                               // (terminated)
		.out_error         (),                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                               // (terminated)
		.out_channel       ()                                                                                    // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (77),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (57),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (58),
		.PKT_TRANS_POSTED          (59),
		.PKT_TRANS_WRITE           (60),
		.PKT_TRANS_READ            (61),
		.PKT_TRANS_LOCK            (62),
		.PKT_SRC_ID_H              (85),
		.PKT_SRC_ID_L              (79),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (86),
		.PKT_BURSTWRAP_H           (69),
		.PKT_BURSTWRAP_L           (67),
		.PKT_BYTE_CNT_H            (66),
		.PKT_BYTE_CNT_L            (64),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (72),
		.PKT_BURST_SIZE_L          (70),
		.ST_CHANNEL_W              (99),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) ch1_yn2_l_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                           //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                //       clk_reset.reset
		.m0_address              (ch1_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ch1_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ch1_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ch1_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ch1_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ch1_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ch1_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ch1_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ch1_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ch1_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ch1_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ch1_yn2_l_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ch1_yn2_l_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ch1_yn2_l_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ch1_yn2_l_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ch1_yn2_l_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src43_ready),                                                    //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src43_valid),                                                    //                .valid
		.cp_data                 (cmd_xbar_demux_001_src43_data),                                                     //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src43_startofpacket),                                            //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src43_endofpacket),                                              //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src43_channel),                                                  //                .channel
		.rf_sink_ready           (ch1_yn2_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ch1_yn2_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ch1_yn2_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ch1_yn2_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ch1_yn2_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ch1_yn2_l_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ch1_yn2_l_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ch1_yn2_l_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ch1_yn2_l_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ch1_yn2_l_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ch1_yn2_l_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ch1_yn2_l_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (ch1_yn2_l_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (ch1_yn2_l_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ch1_yn2_l_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ch1_yn2_l_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                             //     (terminated)
		.m0_writeresponserequest (),                                                                                  //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                               //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ch1_yn2_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                           //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                // clk_reset.reset
		.in_data           (ch1_yn2_l_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ch1_yn2_l_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ch1_yn2_l_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ch1_yn2_l_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ch1_yn2_l_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ch1_yn2_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ch1_yn2_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ch1_yn2_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ch1_yn2_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ch1_yn2_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                             // (terminated)
		.csr_read          (1'b0),                                                                              // (terminated)
		.csr_write         (1'b0),                                                                              // (terminated)
		.csr_readdata      (),                                                                                  // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                              // (terminated)
		.almost_full_data  (),                                                                                  // (terminated)
		.almost_empty_data (),                                                                                  // (terminated)
		.in_empty          (1'b0),                                                                              // (terminated)
		.out_empty         (),                                                                                  // (terminated)
		.in_error          (1'b0),                                                                              // (terminated)
		.out_error         (),                                                                                  // (terminated)
		.in_channel        (1'b0),                                                                              // (terminated)
		.out_channel       ()                                                                                   // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (77),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (57),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (58),
		.PKT_TRANS_POSTED          (59),
		.PKT_TRANS_WRITE           (60),
		.PKT_TRANS_READ            (61),
		.PKT_TRANS_LOCK            (62),
		.PKT_SRC_ID_H              (85),
		.PKT_SRC_ID_L              (79),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (86),
		.PKT_BURSTWRAP_H           (69),
		.PKT_BURSTWRAP_L           (67),
		.PKT_BYTE_CNT_H            (66),
		.PKT_BYTE_CNT_L            (64),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (72),
		.PKT_BURST_SIZE_L          (70),
		.ST_CHANNEL_W              (99),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) ch1_yn3_u_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                           //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                //       clk_reset.reset
		.m0_address              (ch1_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ch1_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ch1_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ch1_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ch1_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ch1_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ch1_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ch1_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ch1_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ch1_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ch1_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ch1_yn3_u_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ch1_yn3_u_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ch1_yn3_u_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ch1_yn3_u_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ch1_yn3_u_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src44_ready),                                                    //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src44_valid),                                                    //                .valid
		.cp_data                 (cmd_xbar_demux_001_src44_data),                                                     //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src44_startofpacket),                                            //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src44_endofpacket),                                              //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src44_channel),                                                  //                .channel
		.rf_sink_ready           (ch1_yn3_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ch1_yn3_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ch1_yn3_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ch1_yn3_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ch1_yn3_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ch1_yn3_u_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ch1_yn3_u_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ch1_yn3_u_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ch1_yn3_u_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ch1_yn3_u_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ch1_yn3_u_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ch1_yn3_u_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (ch1_yn3_u_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (ch1_yn3_u_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ch1_yn3_u_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ch1_yn3_u_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                             //     (terminated)
		.m0_writeresponserequest (),                                                                                  //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                               //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ch1_yn3_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                           //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                // clk_reset.reset
		.in_data           (ch1_yn3_u_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ch1_yn3_u_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ch1_yn3_u_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ch1_yn3_u_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ch1_yn3_u_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ch1_yn3_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ch1_yn3_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ch1_yn3_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ch1_yn3_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ch1_yn3_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                             // (terminated)
		.csr_read          (1'b0),                                                                              // (terminated)
		.csr_write         (1'b0),                                                                              // (terminated)
		.csr_readdata      (),                                                                                  // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                              // (terminated)
		.almost_full_data  (),                                                                                  // (terminated)
		.almost_empty_data (),                                                                                  // (terminated)
		.in_empty          (1'b0),                                                                              // (terminated)
		.out_empty         (),                                                                                  // (terminated)
		.in_error          (1'b0),                                                                              // (terminated)
		.out_error         (),                                                                                  // (terminated)
		.in_channel        (1'b0),                                                                              // (terminated)
		.out_channel       ()                                                                                   // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (77),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (57),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (58),
		.PKT_TRANS_POSTED          (59),
		.PKT_TRANS_WRITE           (60),
		.PKT_TRANS_READ            (61),
		.PKT_TRANS_LOCK            (62),
		.PKT_SRC_ID_H              (85),
		.PKT_SRC_ID_L              (79),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (86),
		.PKT_BURSTWRAP_H           (69),
		.PKT_BURSTWRAP_L           (67),
		.PKT_BYTE_CNT_H            (66),
		.PKT_BYTE_CNT_L            (64),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (72),
		.PKT_BURST_SIZE_L          (70),
		.ST_CHANNEL_W              (99),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) ch1_yn3_mu_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                            //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                 //       clk_reset.reset
		.m0_address              (ch1_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ch1_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ch1_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ch1_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ch1_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ch1_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ch1_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ch1_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ch1_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ch1_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ch1_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ch1_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ch1_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ch1_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ch1_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ch1_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src45_ready),                                                     //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src45_valid),                                                     //                .valid
		.cp_data                 (cmd_xbar_demux_001_src45_data),                                                      //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src45_startofpacket),                                             //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src45_endofpacket),                                               //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src45_channel),                                                   //                .channel
		.rf_sink_ready           (ch1_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ch1_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ch1_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ch1_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ch1_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ch1_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ch1_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ch1_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ch1_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ch1_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ch1_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ch1_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (ch1_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (ch1_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ch1_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ch1_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                              //     (terminated)
		.m0_writeresponserequest (),                                                                                   //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ch1_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                            //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                 // clk_reset.reset
		.in_data           (ch1_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ch1_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ch1_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ch1_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ch1_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ch1_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ch1_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ch1_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ch1_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ch1_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                              // (terminated)
		.csr_read          (1'b0),                                                                               // (terminated)
		.csr_write         (1'b0),                                                                               // (terminated)
		.csr_readdata      (),                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                               // (terminated)
		.almost_full_data  (),                                                                                   // (terminated)
		.almost_empty_data (),                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                               // (terminated)
		.out_empty         (),                                                                                   // (terminated)
		.in_error          (1'b0),                                                                               // (terminated)
		.out_error         (),                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                               // (terminated)
		.out_channel       ()                                                                                    // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (77),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (57),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (58),
		.PKT_TRANS_POSTED          (59),
		.PKT_TRANS_WRITE           (60),
		.PKT_TRANS_READ            (61),
		.PKT_TRANS_LOCK            (62),
		.PKT_SRC_ID_H              (85),
		.PKT_SRC_ID_L              (79),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (86),
		.PKT_BURSTWRAP_H           (69),
		.PKT_BURSTWRAP_L           (67),
		.PKT_BYTE_CNT_H            (66),
		.PKT_BYTE_CNT_L            (64),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (72),
		.PKT_BURST_SIZE_L          (70),
		.ST_CHANNEL_W              (99),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) ch1_yn3_ml_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                            //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                 //       clk_reset.reset
		.m0_address              (ch1_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ch1_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ch1_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ch1_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ch1_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ch1_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ch1_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ch1_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ch1_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ch1_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ch1_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ch1_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ch1_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ch1_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ch1_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ch1_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src46_ready),                                                     //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src46_valid),                                                     //                .valid
		.cp_data                 (cmd_xbar_demux_001_src46_data),                                                      //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src46_startofpacket),                                             //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src46_endofpacket),                                               //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src46_channel),                                                   //                .channel
		.rf_sink_ready           (ch1_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ch1_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ch1_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ch1_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ch1_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ch1_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ch1_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ch1_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ch1_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ch1_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ch1_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ch1_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (ch1_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (ch1_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ch1_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ch1_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                              //     (terminated)
		.m0_writeresponserequest (),                                                                                   //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ch1_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                            //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                 // clk_reset.reset
		.in_data           (ch1_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ch1_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ch1_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ch1_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ch1_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ch1_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ch1_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ch1_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ch1_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ch1_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                              // (terminated)
		.csr_read          (1'b0),                                                                               // (terminated)
		.csr_write         (1'b0),                                                                               // (terminated)
		.csr_readdata      (),                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                               // (terminated)
		.almost_full_data  (),                                                                                   // (terminated)
		.almost_empty_data (),                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                               // (terminated)
		.out_empty         (),                                                                                   // (terminated)
		.in_error          (1'b0),                                                                               // (terminated)
		.out_error         (),                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                               // (terminated)
		.out_channel       ()                                                                                    // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (77),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (57),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (58),
		.PKT_TRANS_POSTED          (59),
		.PKT_TRANS_WRITE           (60),
		.PKT_TRANS_READ            (61),
		.PKT_TRANS_LOCK            (62),
		.PKT_SRC_ID_H              (85),
		.PKT_SRC_ID_L              (79),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (86),
		.PKT_BURSTWRAP_H           (69),
		.PKT_BURSTWRAP_L           (67),
		.PKT_BYTE_CNT_H            (66),
		.PKT_BYTE_CNT_L            (64),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (72),
		.PKT_BURST_SIZE_L          (70),
		.ST_CHANNEL_W              (99),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) ch1_yn3_l_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                           //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                //       clk_reset.reset
		.m0_address              (ch1_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ch1_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ch1_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ch1_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ch1_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ch1_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ch1_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ch1_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ch1_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ch1_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ch1_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ch1_yn3_l_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ch1_yn3_l_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ch1_yn3_l_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ch1_yn3_l_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ch1_yn3_l_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src47_ready),                                                    //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src47_valid),                                                    //                .valid
		.cp_data                 (cmd_xbar_demux_001_src47_data),                                                     //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src47_startofpacket),                                            //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src47_endofpacket),                                              //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src47_channel),                                                  //                .channel
		.rf_sink_ready           (ch1_yn3_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ch1_yn3_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ch1_yn3_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ch1_yn3_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ch1_yn3_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ch1_yn3_l_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ch1_yn3_l_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ch1_yn3_l_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ch1_yn3_l_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ch1_yn3_l_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ch1_yn3_l_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ch1_yn3_l_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (ch1_yn3_l_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (ch1_yn3_l_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ch1_yn3_l_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ch1_yn3_l_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                             //     (terminated)
		.m0_writeresponserequest (),                                                                                  //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                               //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ch1_yn3_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                           //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                // clk_reset.reset
		.in_data           (ch1_yn3_l_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ch1_yn3_l_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ch1_yn3_l_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ch1_yn3_l_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ch1_yn3_l_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ch1_yn3_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ch1_yn3_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ch1_yn3_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ch1_yn3_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ch1_yn3_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                             // (terminated)
		.csr_read          (1'b0),                                                                              // (terminated)
		.csr_write         (1'b0),                                                                              // (terminated)
		.csr_readdata      (),                                                                                  // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                              // (terminated)
		.almost_full_data  (),                                                                                  // (terminated)
		.almost_empty_data (),                                                                                  // (terminated)
		.in_empty          (1'b0),                                                                              // (terminated)
		.out_empty         (),                                                                                  // (terminated)
		.in_error          (1'b0),                                                                              // (terminated)
		.out_error         (),                                                                                  // (terminated)
		.in_channel        (1'b0),                                                                              // (terminated)
		.out_channel       ()                                                                                   // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (77),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (57),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (58),
		.PKT_TRANS_POSTED          (59),
		.PKT_TRANS_WRITE           (60),
		.PKT_TRANS_READ            (61),
		.PKT_TRANS_LOCK            (62),
		.PKT_SRC_ID_H              (85),
		.PKT_SRC_ID_L              (79),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (86),
		.PKT_BURSTWRAP_H           (69),
		.PKT_BURSTWRAP_L           (67),
		.PKT_BYTE_CNT_H            (66),
		.PKT_BYTE_CNT_L            (64),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (72),
		.PKT_BURST_SIZE_L          (70),
		.ST_CHANNEL_W              (99),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) ch2_timer_rst_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                               //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                    //       clk_reset.reset
		.m0_address              (ch2_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ch2_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ch2_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ch2_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ch2_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ch2_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ch2_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ch2_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ch2_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ch2_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ch2_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ch2_timer_rst_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ch2_timer_rst_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ch2_timer_rst_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ch2_timer_rst_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ch2_timer_rst_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src48_ready),                                                        //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src48_valid),                                                        //                .valid
		.cp_data                 (cmd_xbar_demux_001_src48_data),                                                         //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src48_startofpacket),                                                //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src48_endofpacket),                                                  //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src48_channel),                                                      //                .channel
		.rf_sink_ready           (ch2_timer_rst_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ch2_timer_rst_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ch2_timer_rst_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ch2_timer_rst_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ch2_timer_rst_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ch2_timer_rst_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ch2_timer_rst_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ch2_timer_rst_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ch2_timer_rst_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ch2_timer_rst_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ch2_timer_rst_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ch2_timer_rst_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (ch2_timer_rst_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (ch2_timer_rst_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ch2_timer_rst_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ch2_timer_rst_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                 //     (terminated)
		.m0_writeresponserequest (),                                                                                      //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                   //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ch2_timer_rst_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                               //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                    // clk_reset.reset
		.in_data           (ch2_timer_rst_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ch2_timer_rst_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ch2_timer_rst_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ch2_timer_rst_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ch2_timer_rst_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ch2_timer_rst_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ch2_timer_rst_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ch2_timer_rst_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ch2_timer_rst_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ch2_timer_rst_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                 // (terminated)
		.csr_read          (1'b0),                                                                                  // (terminated)
		.csr_write         (1'b0),                                                                                  // (terminated)
		.csr_readdata      (),                                                                                      // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                  // (terminated)
		.almost_full_data  (),                                                                                      // (terminated)
		.almost_empty_data (),                                                                                      // (terminated)
		.in_empty          (1'b0),                                                                                  // (terminated)
		.out_empty         (),                                                                                      // (terminated)
		.in_error          (1'b0),                                                                                  // (terminated)
		.out_error         (),                                                                                      // (terminated)
		.in_channel        (1'b0),                                                                                  // (terminated)
		.out_channel       ()                                                                                       // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (77),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (57),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (58),
		.PKT_TRANS_POSTED          (59),
		.PKT_TRANS_WRITE           (60),
		.PKT_TRANS_READ            (61),
		.PKT_TRANS_LOCK            (62),
		.PKT_SRC_ID_H              (85),
		.PKT_SRC_ID_L              (79),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (86),
		.PKT_BURSTWRAP_H           (69),
		.PKT_BURSTWRAP_L           (67),
		.PKT_BYTE_CNT_H            (66),
		.PKT_BYTE_CNT_L            (64),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (72),
		.PKT_BURST_SIZE_L          (70),
		.ST_CHANNEL_W              (99),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) ch2_thresh_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                            //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                 //       clk_reset.reset
		.m0_address              (ch2_thresh_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ch2_thresh_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ch2_thresh_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ch2_thresh_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ch2_thresh_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ch2_thresh_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ch2_thresh_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ch2_thresh_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ch2_thresh_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ch2_thresh_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ch2_thresh_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ch2_thresh_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ch2_thresh_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ch2_thresh_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ch2_thresh_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ch2_thresh_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src49_ready),                                                     //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src49_valid),                                                     //                .valid
		.cp_data                 (cmd_xbar_demux_001_src49_data),                                                      //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src49_startofpacket),                                             //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src49_endofpacket),                                               //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src49_channel),                                                   //                .channel
		.rf_sink_ready           (ch2_thresh_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ch2_thresh_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ch2_thresh_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ch2_thresh_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ch2_thresh_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ch2_thresh_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ch2_thresh_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ch2_thresh_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ch2_thresh_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ch2_thresh_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ch2_thresh_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ch2_thresh_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (ch2_thresh_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (ch2_thresh_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ch2_thresh_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ch2_thresh_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                              //     (terminated)
		.m0_writeresponserequest (),                                                                                   //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ch2_thresh_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                            //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                 // clk_reset.reset
		.in_data           (ch2_thresh_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ch2_thresh_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ch2_thresh_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ch2_thresh_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ch2_thresh_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ch2_thresh_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ch2_thresh_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ch2_thresh_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ch2_thresh_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ch2_thresh_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                              // (terminated)
		.csr_read          (1'b0),                                                                               // (terminated)
		.csr_write         (1'b0),                                                                               // (terminated)
		.csr_readdata      (),                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                               // (terminated)
		.almost_full_data  (),                                                                                   // (terminated)
		.almost_empty_data (),                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                               // (terminated)
		.out_empty         (),                                                                                   // (terminated)
		.in_error          (1'b0),                                                                               // (terminated)
		.out_error         (),                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                               // (terminated)
		.out_channel       ()                                                                                    // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (77),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (57),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (58),
		.PKT_TRANS_POSTED          (59),
		.PKT_TRANS_WRITE           (60),
		.PKT_TRANS_READ            (61),
		.PKT_TRANS_LOCK            (62),
		.PKT_SRC_ID_H              (85),
		.PKT_SRC_ID_L              (79),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (86),
		.PKT_BURSTWRAP_H           (69),
		.PKT_BURSTWRAP_L           (67),
		.PKT_BYTE_CNT_H            (66),
		.PKT_BYTE_CNT_L            (64),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (72),
		.PKT_BURST_SIZE_L          (70),
		.ST_CHANNEL_W              (99),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) ch2_rd_peak_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                             //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                  //       clk_reset.reset
		.m0_address              (ch2_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ch2_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ch2_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ch2_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ch2_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ch2_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ch2_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ch2_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ch2_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ch2_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ch2_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ch2_rd_peak_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ch2_rd_peak_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ch2_rd_peak_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ch2_rd_peak_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ch2_rd_peak_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src50_ready),                                                      //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src50_valid),                                                      //                .valid
		.cp_data                 (cmd_xbar_demux_001_src50_data),                                                       //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src50_startofpacket),                                              //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src50_endofpacket),                                                //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src50_channel),                                                    //                .channel
		.rf_sink_ready           (ch2_rd_peak_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ch2_rd_peak_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ch2_rd_peak_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ch2_rd_peak_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ch2_rd_peak_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ch2_rd_peak_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ch2_rd_peak_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ch2_rd_peak_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ch2_rd_peak_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ch2_rd_peak_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ch2_rd_peak_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ch2_rd_peak_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (ch2_rd_peak_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (ch2_rd_peak_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ch2_rd_peak_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ch2_rd_peak_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                               //     (terminated)
		.m0_writeresponserequest (),                                                                                    //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                 //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ch2_rd_peak_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                             //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                  // clk_reset.reset
		.in_data           (ch2_rd_peak_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ch2_rd_peak_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ch2_rd_peak_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ch2_rd_peak_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ch2_rd_peak_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ch2_rd_peak_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ch2_rd_peak_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ch2_rd_peak_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ch2_rd_peak_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ch2_rd_peak_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                               // (terminated)
		.csr_read          (1'b0),                                                                                // (terminated)
		.csr_write         (1'b0),                                                                                // (terminated)
		.csr_readdata      (),                                                                                    // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                // (terminated)
		.almost_full_data  (),                                                                                    // (terminated)
		.almost_empty_data (),                                                                                    // (terminated)
		.in_empty          (1'b0),                                                                                // (terminated)
		.out_empty         (),                                                                                    // (terminated)
		.in_error          (1'b0),                                                                                // (terminated)
		.out_error         (),                                                                                    // (terminated)
		.in_channel        (1'b0),                                                                                // (terminated)
		.out_channel       ()                                                                                     // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (77),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (57),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (58),
		.PKT_TRANS_POSTED          (59),
		.PKT_TRANS_WRITE           (60),
		.PKT_TRANS_READ            (61),
		.PKT_TRANS_LOCK            (62),
		.PKT_SRC_ID_H              (85),
		.PKT_SRC_ID_L              (79),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (86),
		.PKT_BURSTWRAP_H           (69),
		.PKT_BURSTWRAP_L           (67),
		.PKT_BYTE_CNT_H            (66),
		.PKT_BYTE_CNT_L            (64),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (72),
		.PKT_BURST_SIZE_L          (70),
		.ST_CHANNEL_W              (99),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) ch2_peak_found_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                     //       clk_reset.reset
		.m0_address              (ch2_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ch2_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ch2_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ch2_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ch2_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ch2_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ch2_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ch2_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ch2_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ch2_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ch2_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ch2_peak_found_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ch2_peak_found_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ch2_peak_found_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ch2_peak_found_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ch2_peak_found_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src51_ready),                                                         //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src51_valid),                                                         //                .valid
		.cp_data                 (cmd_xbar_demux_001_src51_data),                                                          //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src51_startofpacket),                                                 //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src51_endofpacket),                                                   //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src51_channel),                                                       //                .channel
		.rf_sink_ready           (ch2_peak_found_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ch2_peak_found_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ch2_peak_found_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ch2_peak_found_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ch2_peak_found_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ch2_peak_found_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ch2_peak_found_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ch2_peak_found_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ch2_peak_found_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ch2_peak_found_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ch2_peak_found_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ch2_peak_found_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (ch2_peak_found_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (ch2_peak_found_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ch2_peak_found_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ch2_peak_found_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                  //     (terminated)
		.m0_writeresponserequest (),                                                                                       //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                    //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ch2_peak_found_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                     // clk_reset.reset
		.in_data           (ch2_peak_found_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ch2_peak_found_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ch2_peak_found_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ch2_peak_found_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ch2_peak_found_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ch2_peak_found_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ch2_peak_found_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ch2_peak_found_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ch2_peak_found_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ch2_peak_found_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                  // (terminated)
		.csr_read          (1'b0),                                                                                   // (terminated)
		.csr_write         (1'b0),                                                                                   // (terminated)
		.csr_readdata      (),                                                                                       // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                   // (terminated)
		.almost_full_data  (),                                                                                       // (terminated)
		.almost_empty_data (),                                                                                       // (terminated)
		.in_empty          (1'b0),                                                                                   // (terminated)
		.out_empty         (),                                                                                       // (terminated)
		.in_error          (1'b0),                                                                                   // (terminated)
		.out_error         (),                                                                                       // (terminated)
		.in_channel        (1'b0),                                                                                   // (terminated)
		.out_channel       ()                                                                                        // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (77),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (57),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (58),
		.PKT_TRANS_POSTED          (59),
		.PKT_TRANS_WRITE           (60),
		.PKT_TRANS_READ            (61),
		.PKT_TRANS_LOCK            (62),
		.PKT_SRC_ID_H              (85),
		.PKT_SRC_ID_L              (79),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (86),
		.PKT_BURSTWRAP_H           (69),
		.PKT_BURSTWRAP_L           (67),
		.PKT_BYTE_CNT_H            (66),
		.PKT_BYTE_CNT_L            (64),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (72),
		.PKT_BURST_SIZE_L          (70),
		.ST_CHANNEL_W              (99),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) ch2_time_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                          //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                               //       clk_reset.reset
		.m0_address              (ch2_time_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ch2_time_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ch2_time_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ch2_time_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ch2_time_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ch2_time_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ch2_time_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ch2_time_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ch2_time_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ch2_time_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ch2_time_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ch2_time_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ch2_time_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ch2_time_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ch2_time_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ch2_time_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src52_ready),                                                   //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src52_valid),                                                   //                .valid
		.cp_data                 (cmd_xbar_demux_001_src52_data),                                                    //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src52_startofpacket),                                           //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src52_endofpacket),                                             //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src52_channel),                                                 //                .channel
		.rf_sink_ready           (ch2_time_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ch2_time_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ch2_time_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ch2_time_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ch2_time_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ch2_time_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ch2_time_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ch2_time_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ch2_time_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ch2_time_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ch2_time_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ch2_time_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (ch2_time_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (ch2_time_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ch2_time_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ch2_time_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                            //     (terminated)
		.m0_writeresponserequest (),                                                                                 //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                              //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ch2_time_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                          //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                               // clk_reset.reset
		.in_data           (ch2_time_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ch2_time_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ch2_time_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ch2_time_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ch2_time_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ch2_time_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ch2_time_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ch2_time_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ch2_time_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ch2_time_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                            // (terminated)
		.csr_read          (1'b0),                                                                             // (terminated)
		.csr_write         (1'b0),                                                                             // (terminated)
		.csr_readdata      (),                                                                                 // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                             // (terminated)
		.almost_full_data  (),                                                                                 // (terminated)
		.almost_empty_data (),                                                                                 // (terminated)
		.in_empty          (1'b0),                                                                             // (terminated)
		.out_empty         (),                                                                                 // (terminated)
		.in_error          (1'b0),                                                                             // (terminated)
		.out_error         (),                                                                                 // (terminated)
		.in_channel        (1'b0),                                                                             // (terminated)
		.out_channel       ()                                                                                  // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (77),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (57),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (58),
		.PKT_TRANS_POSTED          (59),
		.PKT_TRANS_WRITE           (60),
		.PKT_TRANS_READ            (61),
		.PKT_TRANS_LOCK            (62),
		.PKT_SRC_ID_H              (85),
		.PKT_SRC_ID_L              (79),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (86),
		.PKT_BURSTWRAP_H           (69),
		.PKT_BURSTWRAP_L           (67),
		.PKT_BYTE_CNT_H            (66),
		.PKT_BYTE_CNT_L            (64),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (72),
		.PKT_BURST_SIZE_L          (70),
		.ST_CHANNEL_W              (99),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) ch2_yn1_u_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                           //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                //       clk_reset.reset
		.m0_address              (ch2_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ch2_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ch2_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ch2_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ch2_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ch2_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ch2_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ch2_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ch2_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ch2_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ch2_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ch2_yn1_u_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ch2_yn1_u_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ch2_yn1_u_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ch2_yn1_u_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ch2_yn1_u_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src53_ready),                                                    //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src53_valid),                                                    //                .valid
		.cp_data                 (cmd_xbar_demux_001_src53_data),                                                     //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src53_startofpacket),                                            //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src53_endofpacket),                                              //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src53_channel),                                                  //                .channel
		.rf_sink_ready           (ch2_yn1_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ch2_yn1_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ch2_yn1_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ch2_yn1_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ch2_yn1_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ch2_yn1_u_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ch2_yn1_u_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ch2_yn1_u_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ch2_yn1_u_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ch2_yn1_u_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ch2_yn1_u_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ch2_yn1_u_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (ch2_yn1_u_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (ch2_yn1_u_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ch2_yn1_u_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ch2_yn1_u_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                             //     (terminated)
		.m0_writeresponserequest (),                                                                                  //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                               //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ch2_yn1_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                           //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                // clk_reset.reset
		.in_data           (ch2_yn1_u_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ch2_yn1_u_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ch2_yn1_u_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ch2_yn1_u_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ch2_yn1_u_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ch2_yn1_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ch2_yn1_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ch2_yn1_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ch2_yn1_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ch2_yn1_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                             // (terminated)
		.csr_read          (1'b0),                                                                              // (terminated)
		.csr_write         (1'b0),                                                                              // (terminated)
		.csr_readdata      (),                                                                                  // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                              // (terminated)
		.almost_full_data  (),                                                                                  // (terminated)
		.almost_empty_data (),                                                                                  // (terminated)
		.in_empty          (1'b0),                                                                              // (terminated)
		.out_empty         (),                                                                                  // (terminated)
		.in_error          (1'b0),                                                                              // (terminated)
		.out_error         (),                                                                                  // (terminated)
		.in_channel        (1'b0),                                                                              // (terminated)
		.out_channel       ()                                                                                   // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (77),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (57),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (58),
		.PKT_TRANS_POSTED          (59),
		.PKT_TRANS_WRITE           (60),
		.PKT_TRANS_READ            (61),
		.PKT_TRANS_LOCK            (62),
		.PKT_SRC_ID_H              (85),
		.PKT_SRC_ID_L              (79),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (86),
		.PKT_BURSTWRAP_H           (69),
		.PKT_BURSTWRAP_L           (67),
		.PKT_BYTE_CNT_H            (66),
		.PKT_BYTE_CNT_L            (64),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (72),
		.PKT_BURST_SIZE_L          (70),
		.ST_CHANNEL_W              (99),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) ch2_yn1_mu_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                            //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                 //       clk_reset.reset
		.m0_address              (ch2_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ch2_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ch2_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ch2_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ch2_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ch2_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ch2_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ch2_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ch2_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ch2_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ch2_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ch2_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ch2_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ch2_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ch2_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ch2_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src54_ready),                                                     //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src54_valid),                                                     //                .valid
		.cp_data                 (cmd_xbar_demux_001_src54_data),                                                      //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src54_startofpacket),                                             //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src54_endofpacket),                                               //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src54_channel),                                                   //                .channel
		.rf_sink_ready           (ch2_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ch2_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ch2_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ch2_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ch2_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ch2_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ch2_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ch2_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ch2_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ch2_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ch2_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ch2_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (ch2_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (ch2_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ch2_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ch2_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                              //     (terminated)
		.m0_writeresponserequest (),                                                                                   //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ch2_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                            //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                 // clk_reset.reset
		.in_data           (ch2_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ch2_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ch2_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ch2_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ch2_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ch2_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ch2_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ch2_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ch2_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ch2_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                              // (terminated)
		.csr_read          (1'b0),                                                                               // (terminated)
		.csr_write         (1'b0),                                                                               // (terminated)
		.csr_readdata      (),                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                               // (terminated)
		.almost_full_data  (),                                                                                   // (terminated)
		.almost_empty_data (),                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                               // (terminated)
		.out_empty         (),                                                                                   // (terminated)
		.in_error          (1'b0),                                                                               // (terminated)
		.out_error         (),                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                               // (terminated)
		.out_channel       ()                                                                                    // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (77),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (57),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (58),
		.PKT_TRANS_POSTED          (59),
		.PKT_TRANS_WRITE           (60),
		.PKT_TRANS_READ            (61),
		.PKT_TRANS_LOCK            (62),
		.PKT_SRC_ID_H              (85),
		.PKT_SRC_ID_L              (79),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (86),
		.PKT_BURSTWRAP_H           (69),
		.PKT_BURSTWRAP_L           (67),
		.PKT_BYTE_CNT_H            (66),
		.PKT_BYTE_CNT_L            (64),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (72),
		.PKT_BURST_SIZE_L          (70),
		.ST_CHANNEL_W              (99),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) ch2_yn1_ml_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                            //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                 //       clk_reset.reset
		.m0_address              (ch2_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ch2_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ch2_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ch2_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ch2_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ch2_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ch2_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ch2_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ch2_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ch2_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ch2_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ch2_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ch2_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ch2_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ch2_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ch2_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src55_ready),                                                     //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src55_valid),                                                     //                .valid
		.cp_data                 (cmd_xbar_demux_001_src55_data),                                                      //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src55_startofpacket),                                             //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src55_endofpacket),                                               //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src55_channel),                                                   //                .channel
		.rf_sink_ready           (ch2_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ch2_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ch2_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ch2_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ch2_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ch2_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ch2_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ch2_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ch2_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ch2_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ch2_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ch2_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (ch2_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (ch2_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ch2_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ch2_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                              //     (terminated)
		.m0_writeresponserequest (),                                                                                   //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ch2_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                            //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                 // clk_reset.reset
		.in_data           (ch2_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ch2_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ch2_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ch2_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ch2_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ch2_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ch2_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ch2_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ch2_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ch2_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                              // (terminated)
		.csr_read          (1'b0),                                                                               // (terminated)
		.csr_write         (1'b0),                                                                               // (terminated)
		.csr_readdata      (),                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                               // (terminated)
		.almost_full_data  (),                                                                                   // (terminated)
		.almost_empty_data (),                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                               // (terminated)
		.out_empty         (),                                                                                   // (terminated)
		.in_error          (1'b0),                                                                               // (terminated)
		.out_error         (),                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                               // (terminated)
		.out_channel       ()                                                                                    // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (77),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (57),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (58),
		.PKT_TRANS_POSTED          (59),
		.PKT_TRANS_WRITE           (60),
		.PKT_TRANS_READ            (61),
		.PKT_TRANS_LOCK            (62),
		.PKT_SRC_ID_H              (85),
		.PKT_SRC_ID_L              (79),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (86),
		.PKT_BURSTWRAP_H           (69),
		.PKT_BURSTWRAP_L           (67),
		.PKT_BYTE_CNT_H            (66),
		.PKT_BYTE_CNT_L            (64),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (72),
		.PKT_BURST_SIZE_L          (70),
		.ST_CHANNEL_W              (99),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) ch2_yn1_l_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                           //             clk.clk
		.reset                   (nios_cpu_jtag_debug_module_reset_reset),                                            //       clk_reset.reset
		.m0_address              (ch2_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ch2_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ch2_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ch2_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ch2_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ch2_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ch2_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ch2_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ch2_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ch2_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ch2_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ch2_yn1_l_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ch2_yn1_l_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ch2_yn1_l_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ch2_yn1_l_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ch2_yn1_l_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src56_ready),                                                    //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src56_valid),                                                    //                .valid
		.cp_data                 (cmd_xbar_demux_001_src56_data),                                                     //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src56_startofpacket),                                            //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src56_endofpacket),                                              //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src56_channel),                                                  //                .channel
		.rf_sink_ready           (ch2_yn1_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ch2_yn1_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ch2_yn1_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ch2_yn1_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ch2_yn1_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ch2_yn1_l_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ch2_yn1_l_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ch2_yn1_l_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ch2_yn1_l_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ch2_yn1_l_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ch2_yn1_l_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ch2_yn1_l_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (ch2_yn1_l_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (ch2_yn1_l_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ch2_yn1_l_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ch2_yn1_l_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                             //     (terminated)
		.m0_writeresponserequest (),                                                                                  //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                               //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ch2_yn1_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                           //       clk.clk
		.reset             (nios_cpu_jtag_debug_module_reset_reset),                                            // clk_reset.reset
		.in_data           (ch2_yn1_l_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ch2_yn1_l_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ch2_yn1_l_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ch2_yn1_l_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ch2_yn1_l_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ch2_yn1_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ch2_yn1_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ch2_yn1_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ch2_yn1_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ch2_yn1_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                             // (terminated)
		.csr_read          (1'b0),                                                                              // (terminated)
		.csr_write         (1'b0),                                                                              // (terminated)
		.csr_readdata      (),                                                                                  // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                              // (terminated)
		.almost_full_data  (),                                                                                  // (terminated)
		.almost_empty_data (),                                                                                  // (terminated)
		.in_empty          (1'b0),                                                                              // (terminated)
		.out_empty         (),                                                                                  // (terminated)
		.in_error          (1'b0),                                                                              // (terminated)
		.out_error         (),                                                                                  // (terminated)
		.in_channel        (1'b0),                                                                              // (terminated)
		.out_channel       ()                                                                                   // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (77),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (57),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (58),
		.PKT_TRANS_POSTED          (59),
		.PKT_TRANS_WRITE           (60),
		.PKT_TRANS_READ            (61),
		.PKT_TRANS_LOCK            (62),
		.PKT_SRC_ID_H              (85),
		.PKT_SRC_ID_L              (79),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (86),
		.PKT_BURSTWRAP_H           (69),
		.PKT_BURSTWRAP_L           (67),
		.PKT_BYTE_CNT_H            (66),
		.PKT_BYTE_CNT_L            (64),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (72),
		.PKT_BURST_SIZE_L          (70),
		.ST_CHANNEL_W              (99),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) ch2_yn2_u_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                           //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                //       clk_reset.reset
		.m0_address              (ch2_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ch2_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ch2_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ch2_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ch2_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ch2_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ch2_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ch2_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ch2_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ch2_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ch2_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ch2_yn2_u_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ch2_yn2_u_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ch2_yn2_u_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ch2_yn2_u_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ch2_yn2_u_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src57_ready),                                                    //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src57_valid),                                                    //                .valid
		.cp_data                 (cmd_xbar_demux_001_src57_data),                                                     //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src57_startofpacket),                                            //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src57_endofpacket),                                              //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src57_channel),                                                  //                .channel
		.rf_sink_ready           (ch2_yn2_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ch2_yn2_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ch2_yn2_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ch2_yn2_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ch2_yn2_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ch2_yn2_u_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ch2_yn2_u_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ch2_yn2_u_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ch2_yn2_u_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ch2_yn2_u_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ch2_yn2_u_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ch2_yn2_u_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (ch2_yn2_u_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (ch2_yn2_u_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ch2_yn2_u_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ch2_yn2_u_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                             //     (terminated)
		.m0_writeresponserequest (),                                                                                  //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                               //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ch2_yn2_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                           //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                // clk_reset.reset
		.in_data           (ch2_yn2_u_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ch2_yn2_u_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ch2_yn2_u_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ch2_yn2_u_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ch2_yn2_u_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ch2_yn2_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ch2_yn2_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ch2_yn2_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ch2_yn2_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ch2_yn2_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                             // (terminated)
		.csr_read          (1'b0),                                                                              // (terminated)
		.csr_write         (1'b0),                                                                              // (terminated)
		.csr_readdata      (),                                                                                  // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                              // (terminated)
		.almost_full_data  (),                                                                                  // (terminated)
		.almost_empty_data (),                                                                                  // (terminated)
		.in_empty          (1'b0),                                                                              // (terminated)
		.out_empty         (),                                                                                  // (terminated)
		.in_error          (1'b0),                                                                              // (terminated)
		.out_error         (),                                                                                  // (terminated)
		.in_channel        (1'b0),                                                                              // (terminated)
		.out_channel       ()                                                                                   // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (77),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (57),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (58),
		.PKT_TRANS_POSTED          (59),
		.PKT_TRANS_WRITE           (60),
		.PKT_TRANS_READ            (61),
		.PKT_TRANS_LOCK            (62),
		.PKT_SRC_ID_H              (85),
		.PKT_SRC_ID_L              (79),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (86),
		.PKT_BURSTWRAP_H           (69),
		.PKT_BURSTWRAP_L           (67),
		.PKT_BYTE_CNT_H            (66),
		.PKT_BYTE_CNT_L            (64),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (72),
		.PKT_BURST_SIZE_L          (70),
		.ST_CHANNEL_W              (99),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) ch2_yn2_mu_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                            //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                 //       clk_reset.reset
		.m0_address              (ch2_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ch2_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ch2_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ch2_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ch2_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ch2_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ch2_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ch2_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ch2_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ch2_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ch2_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ch2_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ch2_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ch2_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ch2_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ch2_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src58_ready),                                                     //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src58_valid),                                                     //                .valid
		.cp_data                 (cmd_xbar_demux_001_src58_data),                                                      //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src58_startofpacket),                                             //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src58_endofpacket),                                               //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src58_channel),                                                   //                .channel
		.rf_sink_ready           (ch2_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ch2_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ch2_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ch2_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ch2_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ch2_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ch2_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ch2_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ch2_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ch2_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ch2_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ch2_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (ch2_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (ch2_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ch2_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ch2_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                              //     (terminated)
		.m0_writeresponserequest (),                                                                                   //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ch2_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                            //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                 // clk_reset.reset
		.in_data           (ch2_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ch2_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ch2_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ch2_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ch2_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ch2_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ch2_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ch2_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ch2_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ch2_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                              // (terminated)
		.csr_read          (1'b0),                                                                               // (terminated)
		.csr_write         (1'b0),                                                                               // (terminated)
		.csr_readdata      (),                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                               // (terminated)
		.almost_full_data  (),                                                                                   // (terminated)
		.almost_empty_data (),                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                               // (terminated)
		.out_empty         (),                                                                                   // (terminated)
		.in_error          (1'b0),                                                                               // (terminated)
		.out_error         (),                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                               // (terminated)
		.out_channel       ()                                                                                    // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (77),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (57),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (58),
		.PKT_TRANS_POSTED          (59),
		.PKT_TRANS_WRITE           (60),
		.PKT_TRANS_READ            (61),
		.PKT_TRANS_LOCK            (62),
		.PKT_SRC_ID_H              (85),
		.PKT_SRC_ID_L              (79),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (86),
		.PKT_BURSTWRAP_H           (69),
		.PKT_BURSTWRAP_L           (67),
		.PKT_BYTE_CNT_H            (66),
		.PKT_BYTE_CNT_L            (64),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (72),
		.PKT_BURST_SIZE_L          (70),
		.ST_CHANNEL_W              (99),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) ch2_yn2_ml_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                            //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                 //       clk_reset.reset
		.m0_address              (ch2_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ch2_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ch2_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ch2_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ch2_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ch2_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ch2_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ch2_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ch2_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ch2_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ch2_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ch2_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ch2_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ch2_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ch2_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ch2_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src59_ready),                                                     //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src59_valid),                                                     //                .valid
		.cp_data                 (cmd_xbar_demux_001_src59_data),                                                      //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src59_startofpacket),                                             //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src59_endofpacket),                                               //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src59_channel),                                                   //                .channel
		.rf_sink_ready           (ch2_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ch2_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ch2_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ch2_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ch2_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ch2_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ch2_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ch2_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ch2_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ch2_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ch2_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ch2_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (ch2_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (ch2_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ch2_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ch2_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                              //     (terminated)
		.m0_writeresponserequest (),                                                                                   //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ch2_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                            //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                 // clk_reset.reset
		.in_data           (ch2_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ch2_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ch2_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ch2_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ch2_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ch2_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ch2_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ch2_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ch2_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ch2_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                              // (terminated)
		.csr_read          (1'b0),                                                                               // (terminated)
		.csr_write         (1'b0),                                                                               // (terminated)
		.csr_readdata      (),                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                               // (terminated)
		.almost_full_data  (),                                                                                   // (terminated)
		.almost_empty_data (),                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                               // (terminated)
		.out_empty         (),                                                                                   // (terminated)
		.in_error          (1'b0),                                                                               // (terminated)
		.out_error         (),                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                               // (terminated)
		.out_channel       ()                                                                                    // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (77),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (57),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (58),
		.PKT_TRANS_POSTED          (59),
		.PKT_TRANS_WRITE           (60),
		.PKT_TRANS_READ            (61),
		.PKT_TRANS_LOCK            (62),
		.PKT_SRC_ID_H              (85),
		.PKT_SRC_ID_L              (79),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (86),
		.PKT_BURSTWRAP_H           (69),
		.PKT_BURSTWRAP_L           (67),
		.PKT_BYTE_CNT_H            (66),
		.PKT_BYTE_CNT_L            (64),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (72),
		.PKT_BURST_SIZE_L          (70),
		.ST_CHANNEL_W              (99),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) ch2_yn2_l_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                           //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                //       clk_reset.reset
		.m0_address              (ch2_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ch2_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ch2_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ch2_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ch2_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ch2_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ch2_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ch2_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ch2_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ch2_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ch2_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ch2_yn2_l_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ch2_yn2_l_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ch2_yn2_l_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ch2_yn2_l_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ch2_yn2_l_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src60_ready),                                                    //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src60_valid),                                                    //                .valid
		.cp_data                 (cmd_xbar_demux_001_src60_data),                                                     //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src60_startofpacket),                                            //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src60_endofpacket),                                              //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src60_channel),                                                  //                .channel
		.rf_sink_ready           (ch2_yn2_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ch2_yn2_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ch2_yn2_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ch2_yn2_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ch2_yn2_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ch2_yn2_l_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ch2_yn2_l_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ch2_yn2_l_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ch2_yn2_l_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ch2_yn2_l_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ch2_yn2_l_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ch2_yn2_l_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (ch2_yn2_l_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (ch2_yn2_l_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ch2_yn2_l_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ch2_yn2_l_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                             //     (terminated)
		.m0_writeresponserequest (),                                                                                  //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                               //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ch2_yn2_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                           //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                // clk_reset.reset
		.in_data           (ch2_yn2_l_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ch2_yn2_l_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ch2_yn2_l_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ch2_yn2_l_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ch2_yn2_l_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ch2_yn2_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ch2_yn2_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ch2_yn2_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ch2_yn2_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ch2_yn2_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                             // (terminated)
		.csr_read          (1'b0),                                                                              // (terminated)
		.csr_write         (1'b0),                                                                              // (terminated)
		.csr_readdata      (),                                                                                  // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                              // (terminated)
		.almost_full_data  (),                                                                                  // (terminated)
		.almost_empty_data (),                                                                                  // (terminated)
		.in_empty          (1'b0),                                                                              // (terminated)
		.out_empty         (),                                                                                  // (terminated)
		.in_error          (1'b0),                                                                              // (terminated)
		.out_error         (),                                                                                  // (terminated)
		.in_channel        (1'b0),                                                                              // (terminated)
		.out_channel       ()                                                                                   // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (77),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (57),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (58),
		.PKT_TRANS_POSTED          (59),
		.PKT_TRANS_WRITE           (60),
		.PKT_TRANS_READ            (61),
		.PKT_TRANS_LOCK            (62),
		.PKT_SRC_ID_H              (85),
		.PKT_SRC_ID_L              (79),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (86),
		.PKT_BURSTWRAP_H           (69),
		.PKT_BURSTWRAP_L           (67),
		.PKT_BYTE_CNT_H            (66),
		.PKT_BYTE_CNT_L            (64),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (72),
		.PKT_BURST_SIZE_L          (70),
		.ST_CHANNEL_W              (99),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) ch2_yn3_u_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                           //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                //       clk_reset.reset
		.m0_address              (ch2_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ch2_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ch2_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ch2_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ch2_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ch2_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ch2_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ch2_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ch2_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ch2_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ch2_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ch2_yn3_u_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ch2_yn3_u_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ch2_yn3_u_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ch2_yn3_u_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ch2_yn3_u_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src61_ready),                                                    //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src61_valid),                                                    //                .valid
		.cp_data                 (cmd_xbar_demux_001_src61_data),                                                     //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src61_startofpacket),                                            //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src61_endofpacket),                                              //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src61_channel),                                                  //                .channel
		.rf_sink_ready           (ch2_yn3_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ch2_yn3_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ch2_yn3_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ch2_yn3_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ch2_yn3_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ch2_yn3_u_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ch2_yn3_u_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ch2_yn3_u_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ch2_yn3_u_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ch2_yn3_u_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ch2_yn3_u_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ch2_yn3_u_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (ch2_yn3_u_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (ch2_yn3_u_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ch2_yn3_u_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ch2_yn3_u_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                             //     (terminated)
		.m0_writeresponserequest (),                                                                                  //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                               //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ch2_yn3_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                           //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                // clk_reset.reset
		.in_data           (ch2_yn3_u_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ch2_yn3_u_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ch2_yn3_u_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ch2_yn3_u_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ch2_yn3_u_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ch2_yn3_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ch2_yn3_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ch2_yn3_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ch2_yn3_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ch2_yn3_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                             // (terminated)
		.csr_read          (1'b0),                                                                              // (terminated)
		.csr_write         (1'b0),                                                                              // (terminated)
		.csr_readdata      (),                                                                                  // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                              // (terminated)
		.almost_full_data  (),                                                                                  // (terminated)
		.almost_empty_data (),                                                                                  // (terminated)
		.in_empty          (1'b0),                                                                              // (terminated)
		.out_empty         (),                                                                                  // (terminated)
		.in_error          (1'b0),                                                                              // (terminated)
		.out_error         (),                                                                                  // (terminated)
		.in_channel        (1'b0),                                                                              // (terminated)
		.out_channel       ()                                                                                   // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (77),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (57),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (58),
		.PKT_TRANS_POSTED          (59),
		.PKT_TRANS_WRITE           (60),
		.PKT_TRANS_READ            (61),
		.PKT_TRANS_LOCK            (62),
		.PKT_SRC_ID_H              (85),
		.PKT_SRC_ID_L              (79),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (86),
		.PKT_BURSTWRAP_H           (69),
		.PKT_BURSTWRAP_L           (67),
		.PKT_BYTE_CNT_H            (66),
		.PKT_BYTE_CNT_L            (64),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (72),
		.PKT_BURST_SIZE_L          (70),
		.ST_CHANNEL_W              (99),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) ch2_yn3_mu_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                            //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                 //       clk_reset.reset
		.m0_address              (ch2_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ch2_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ch2_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ch2_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ch2_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ch2_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ch2_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ch2_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ch2_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ch2_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ch2_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ch2_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ch2_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ch2_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ch2_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ch2_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src62_ready),                                                     //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src62_valid),                                                     //                .valid
		.cp_data                 (cmd_xbar_demux_001_src62_data),                                                      //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src62_startofpacket),                                             //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src62_endofpacket),                                               //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src62_channel),                                                   //                .channel
		.rf_sink_ready           (ch2_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ch2_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ch2_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ch2_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ch2_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ch2_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ch2_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ch2_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ch2_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ch2_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ch2_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ch2_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (ch2_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (ch2_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ch2_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ch2_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                              //     (terminated)
		.m0_writeresponserequest (),                                                                                   //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ch2_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                            //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                 // clk_reset.reset
		.in_data           (ch2_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ch2_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ch2_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ch2_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ch2_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ch2_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ch2_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ch2_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ch2_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ch2_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                              // (terminated)
		.csr_read          (1'b0),                                                                               // (terminated)
		.csr_write         (1'b0),                                                                               // (terminated)
		.csr_readdata      (),                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                               // (terminated)
		.almost_full_data  (),                                                                                   // (terminated)
		.almost_empty_data (),                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                               // (terminated)
		.out_empty         (),                                                                                   // (terminated)
		.in_error          (1'b0),                                                                               // (terminated)
		.out_error         (),                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                               // (terminated)
		.out_channel       ()                                                                                    // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (77),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (57),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (58),
		.PKT_TRANS_POSTED          (59),
		.PKT_TRANS_WRITE           (60),
		.PKT_TRANS_READ            (61),
		.PKT_TRANS_LOCK            (62),
		.PKT_SRC_ID_H              (85),
		.PKT_SRC_ID_L              (79),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (86),
		.PKT_BURSTWRAP_H           (69),
		.PKT_BURSTWRAP_L           (67),
		.PKT_BYTE_CNT_H            (66),
		.PKT_BYTE_CNT_L            (64),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (72),
		.PKT_BURST_SIZE_L          (70),
		.ST_CHANNEL_W              (99),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) ch2_yn3_ml_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                            //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                 //       clk_reset.reset
		.m0_address              (ch2_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ch2_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ch2_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ch2_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ch2_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ch2_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ch2_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ch2_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ch2_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ch2_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ch2_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ch2_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ch2_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ch2_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ch2_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ch2_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src63_ready),                                                     //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src63_valid),                                                     //                .valid
		.cp_data                 (cmd_xbar_demux_001_src63_data),                                                      //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src63_startofpacket),                                             //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src63_endofpacket),                                               //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src63_channel),                                                   //                .channel
		.rf_sink_ready           (ch2_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ch2_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ch2_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ch2_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ch2_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ch2_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ch2_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ch2_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ch2_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ch2_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ch2_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ch2_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (ch2_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (ch2_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ch2_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ch2_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                              //     (terminated)
		.m0_writeresponserequest (),                                                                                   //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ch2_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                            //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                 // clk_reset.reset
		.in_data           (ch2_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ch2_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ch2_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ch2_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ch2_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ch2_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ch2_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ch2_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ch2_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ch2_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                              // (terminated)
		.csr_read          (1'b0),                                                                               // (terminated)
		.csr_write         (1'b0),                                                                               // (terminated)
		.csr_readdata      (),                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                               // (terminated)
		.almost_full_data  (),                                                                                   // (terminated)
		.almost_empty_data (),                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                               // (terminated)
		.out_empty         (),                                                                                   // (terminated)
		.in_error          (1'b0),                                                                               // (terminated)
		.out_error         (),                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                               // (terminated)
		.out_channel       ()                                                                                    // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (77),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (57),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (58),
		.PKT_TRANS_POSTED          (59),
		.PKT_TRANS_WRITE           (60),
		.PKT_TRANS_READ            (61),
		.PKT_TRANS_LOCK            (62),
		.PKT_SRC_ID_H              (85),
		.PKT_SRC_ID_L              (79),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (86),
		.PKT_BURSTWRAP_H           (69),
		.PKT_BURSTWRAP_L           (67),
		.PKT_BYTE_CNT_H            (66),
		.PKT_BYTE_CNT_L            (64),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (72),
		.PKT_BURST_SIZE_L          (70),
		.ST_CHANNEL_W              (99),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) ch2_yn3_l_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                           //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                //       clk_reset.reset
		.m0_address              (ch2_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ch2_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ch2_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ch2_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ch2_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ch2_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ch2_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ch2_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ch2_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ch2_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ch2_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ch2_yn3_l_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ch2_yn3_l_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ch2_yn3_l_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ch2_yn3_l_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ch2_yn3_l_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src64_ready),                                                    //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src64_valid),                                                    //                .valid
		.cp_data                 (cmd_xbar_demux_001_src64_data),                                                     //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src64_startofpacket),                                            //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src64_endofpacket),                                              //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src64_channel),                                                  //                .channel
		.rf_sink_ready           (ch2_yn3_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ch2_yn3_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ch2_yn3_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ch2_yn3_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ch2_yn3_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ch2_yn3_l_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ch2_yn3_l_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ch2_yn3_l_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ch2_yn3_l_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ch2_yn3_l_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ch2_yn3_l_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ch2_yn3_l_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (ch2_yn3_l_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (ch2_yn3_l_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ch2_yn3_l_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ch2_yn3_l_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                             //     (terminated)
		.m0_writeresponserequest (),                                                                                  //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                               //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ch2_yn3_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                           //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                // clk_reset.reset
		.in_data           (ch2_yn3_l_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ch2_yn3_l_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ch2_yn3_l_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ch2_yn3_l_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ch2_yn3_l_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ch2_yn3_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ch2_yn3_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ch2_yn3_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ch2_yn3_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ch2_yn3_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                             // (terminated)
		.csr_read          (1'b0),                                                                              // (terminated)
		.csr_write         (1'b0),                                                                              // (terminated)
		.csr_readdata      (),                                                                                  // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                              // (terminated)
		.almost_full_data  (),                                                                                  // (terminated)
		.almost_empty_data (),                                                                                  // (terminated)
		.in_empty          (1'b0),                                                                              // (terminated)
		.out_empty         (),                                                                                  // (terminated)
		.in_error          (1'b0),                                                                              // (terminated)
		.out_error         (),                                                                                  // (terminated)
		.in_channel        (1'b0),                                                                              // (terminated)
		.out_channel       ()                                                                                   // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (77),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (57),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (58),
		.PKT_TRANS_POSTED          (59),
		.PKT_TRANS_WRITE           (60),
		.PKT_TRANS_READ            (61),
		.PKT_TRANS_LOCK            (62),
		.PKT_SRC_ID_H              (85),
		.PKT_SRC_ID_L              (79),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (86),
		.PKT_BURSTWRAP_H           (69),
		.PKT_BURSTWRAP_L           (67),
		.PKT_BYTE_CNT_H            (66),
		.PKT_BYTE_CNT_L            (64),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (72),
		.PKT_BURST_SIZE_L          (70),
		.ST_CHANNEL_W              (99),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) ch3_timer_rst_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                               //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                    //       clk_reset.reset
		.m0_address              (ch3_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ch3_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ch3_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ch3_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ch3_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ch3_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ch3_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ch3_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ch3_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ch3_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ch3_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ch3_timer_rst_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ch3_timer_rst_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ch3_timer_rst_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ch3_timer_rst_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ch3_timer_rst_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src65_ready),                                                        //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src65_valid),                                                        //                .valid
		.cp_data                 (cmd_xbar_demux_001_src65_data),                                                         //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src65_startofpacket),                                                //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src65_endofpacket),                                                  //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src65_channel),                                                      //                .channel
		.rf_sink_ready           (ch3_timer_rst_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ch3_timer_rst_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ch3_timer_rst_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ch3_timer_rst_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ch3_timer_rst_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ch3_timer_rst_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ch3_timer_rst_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ch3_timer_rst_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ch3_timer_rst_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ch3_timer_rst_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ch3_timer_rst_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ch3_timer_rst_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (ch3_timer_rst_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (ch3_timer_rst_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ch3_timer_rst_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ch3_timer_rst_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                 //     (terminated)
		.m0_writeresponserequest (),                                                                                      //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                   //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ch3_timer_rst_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                               //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                    // clk_reset.reset
		.in_data           (ch3_timer_rst_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ch3_timer_rst_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ch3_timer_rst_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ch3_timer_rst_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ch3_timer_rst_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ch3_timer_rst_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ch3_timer_rst_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ch3_timer_rst_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ch3_timer_rst_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ch3_timer_rst_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                 // (terminated)
		.csr_read          (1'b0),                                                                                  // (terminated)
		.csr_write         (1'b0),                                                                                  // (terminated)
		.csr_readdata      (),                                                                                      // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                  // (terminated)
		.almost_full_data  (),                                                                                      // (terminated)
		.almost_empty_data (),                                                                                      // (terminated)
		.in_empty          (1'b0),                                                                                  // (terminated)
		.out_empty         (),                                                                                      // (terminated)
		.in_error          (1'b0),                                                                                  // (terminated)
		.out_error         (),                                                                                      // (terminated)
		.in_channel        (1'b0),                                                                                  // (terminated)
		.out_channel       ()                                                                                       // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (77),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (57),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (58),
		.PKT_TRANS_POSTED          (59),
		.PKT_TRANS_WRITE           (60),
		.PKT_TRANS_READ            (61),
		.PKT_TRANS_LOCK            (62),
		.PKT_SRC_ID_H              (85),
		.PKT_SRC_ID_L              (79),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (86),
		.PKT_BURSTWRAP_H           (69),
		.PKT_BURSTWRAP_L           (67),
		.PKT_BYTE_CNT_H            (66),
		.PKT_BYTE_CNT_L            (64),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (72),
		.PKT_BURST_SIZE_L          (70),
		.ST_CHANNEL_W              (99),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) ch3_thresh_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                            //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                 //       clk_reset.reset
		.m0_address              (ch3_thresh_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ch3_thresh_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ch3_thresh_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ch3_thresh_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ch3_thresh_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ch3_thresh_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ch3_thresh_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ch3_thresh_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ch3_thresh_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ch3_thresh_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ch3_thresh_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ch3_thresh_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ch3_thresh_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ch3_thresh_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ch3_thresh_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ch3_thresh_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src66_ready),                                                     //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src66_valid),                                                     //                .valid
		.cp_data                 (cmd_xbar_demux_001_src66_data),                                                      //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src66_startofpacket),                                             //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src66_endofpacket),                                               //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src66_channel),                                                   //                .channel
		.rf_sink_ready           (ch3_thresh_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ch3_thresh_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ch3_thresh_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ch3_thresh_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ch3_thresh_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ch3_thresh_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ch3_thresh_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ch3_thresh_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ch3_thresh_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ch3_thresh_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ch3_thresh_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ch3_thresh_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (ch3_thresh_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (ch3_thresh_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ch3_thresh_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ch3_thresh_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                              //     (terminated)
		.m0_writeresponserequest (),                                                                                   //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ch3_thresh_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                            //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                 // clk_reset.reset
		.in_data           (ch3_thresh_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ch3_thresh_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ch3_thresh_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ch3_thresh_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ch3_thresh_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ch3_thresh_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ch3_thresh_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ch3_thresh_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ch3_thresh_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ch3_thresh_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                              // (terminated)
		.csr_read          (1'b0),                                                                               // (terminated)
		.csr_write         (1'b0),                                                                               // (terminated)
		.csr_readdata      (),                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                               // (terminated)
		.almost_full_data  (),                                                                                   // (terminated)
		.almost_empty_data (),                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                               // (terminated)
		.out_empty         (),                                                                                   // (terminated)
		.in_error          (1'b0),                                                                               // (terminated)
		.out_error         (),                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                               // (terminated)
		.out_channel       ()                                                                                    // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (77),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (57),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (58),
		.PKT_TRANS_POSTED          (59),
		.PKT_TRANS_WRITE           (60),
		.PKT_TRANS_READ            (61),
		.PKT_TRANS_LOCK            (62),
		.PKT_SRC_ID_H              (85),
		.PKT_SRC_ID_L              (79),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (86),
		.PKT_BURSTWRAP_H           (69),
		.PKT_BURSTWRAP_L           (67),
		.PKT_BYTE_CNT_H            (66),
		.PKT_BYTE_CNT_L            (64),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (72),
		.PKT_BURST_SIZE_L          (70),
		.ST_CHANNEL_W              (99),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) ch3_rd_peak_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                             //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                  //       clk_reset.reset
		.m0_address              (ch3_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ch3_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ch3_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ch3_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ch3_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ch3_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ch3_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ch3_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ch3_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ch3_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ch3_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ch3_rd_peak_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ch3_rd_peak_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ch3_rd_peak_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ch3_rd_peak_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ch3_rd_peak_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src67_ready),                                                      //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src67_valid),                                                      //                .valid
		.cp_data                 (cmd_xbar_demux_001_src67_data),                                                       //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src67_startofpacket),                                              //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src67_endofpacket),                                                //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src67_channel),                                                    //                .channel
		.rf_sink_ready           (ch3_rd_peak_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ch3_rd_peak_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ch3_rd_peak_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ch3_rd_peak_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ch3_rd_peak_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ch3_rd_peak_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ch3_rd_peak_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ch3_rd_peak_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ch3_rd_peak_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ch3_rd_peak_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ch3_rd_peak_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ch3_rd_peak_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (ch3_rd_peak_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (ch3_rd_peak_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ch3_rd_peak_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ch3_rd_peak_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                               //     (terminated)
		.m0_writeresponserequest (),                                                                                    //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                 //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ch3_rd_peak_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                             //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                  // clk_reset.reset
		.in_data           (ch3_rd_peak_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ch3_rd_peak_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ch3_rd_peak_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ch3_rd_peak_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ch3_rd_peak_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ch3_rd_peak_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ch3_rd_peak_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ch3_rd_peak_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ch3_rd_peak_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ch3_rd_peak_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                               // (terminated)
		.csr_read          (1'b0),                                                                                // (terminated)
		.csr_write         (1'b0),                                                                                // (terminated)
		.csr_readdata      (),                                                                                    // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                // (terminated)
		.almost_full_data  (),                                                                                    // (terminated)
		.almost_empty_data (),                                                                                    // (terminated)
		.in_empty          (1'b0),                                                                                // (terminated)
		.out_empty         (),                                                                                    // (terminated)
		.in_error          (1'b0),                                                                                // (terminated)
		.out_error         (),                                                                                    // (terminated)
		.in_channel        (1'b0),                                                                                // (terminated)
		.out_channel       ()                                                                                     // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (77),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (57),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (58),
		.PKT_TRANS_POSTED          (59),
		.PKT_TRANS_WRITE           (60),
		.PKT_TRANS_READ            (61),
		.PKT_TRANS_LOCK            (62),
		.PKT_SRC_ID_H              (85),
		.PKT_SRC_ID_L              (79),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (86),
		.PKT_BURSTWRAP_H           (69),
		.PKT_BURSTWRAP_L           (67),
		.PKT_BYTE_CNT_H            (66),
		.PKT_BYTE_CNT_L            (64),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (72),
		.PKT_BURST_SIZE_L          (70),
		.ST_CHANNEL_W              (99),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) ch3_peak_found_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                     //       clk_reset.reset
		.m0_address              (ch3_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ch3_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ch3_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ch3_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ch3_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ch3_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ch3_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ch3_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ch3_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ch3_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ch3_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ch3_peak_found_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ch3_peak_found_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ch3_peak_found_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ch3_peak_found_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ch3_peak_found_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src68_ready),                                                         //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src68_valid),                                                         //                .valid
		.cp_data                 (cmd_xbar_demux_001_src68_data),                                                          //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src68_startofpacket),                                                 //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src68_endofpacket),                                                   //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src68_channel),                                                       //                .channel
		.rf_sink_ready           (ch3_peak_found_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ch3_peak_found_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ch3_peak_found_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ch3_peak_found_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ch3_peak_found_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ch3_peak_found_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ch3_peak_found_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ch3_peak_found_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ch3_peak_found_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ch3_peak_found_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ch3_peak_found_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ch3_peak_found_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (ch3_peak_found_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (ch3_peak_found_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ch3_peak_found_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ch3_peak_found_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                  //     (terminated)
		.m0_writeresponserequest (),                                                                                       //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                    //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ch3_peak_found_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                     // clk_reset.reset
		.in_data           (ch3_peak_found_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ch3_peak_found_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ch3_peak_found_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ch3_peak_found_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ch3_peak_found_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ch3_peak_found_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ch3_peak_found_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ch3_peak_found_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ch3_peak_found_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ch3_peak_found_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                  // (terminated)
		.csr_read          (1'b0),                                                                                   // (terminated)
		.csr_write         (1'b0),                                                                                   // (terminated)
		.csr_readdata      (),                                                                                       // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                   // (terminated)
		.almost_full_data  (),                                                                                       // (terminated)
		.almost_empty_data (),                                                                                       // (terminated)
		.in_empty          (1'b0),                                                                                   // (terminated)
		.out_empty         (),                                                                                       // (terminated)
		.in_error          (1'b0),                                                                                   // (terminated)
		.out_error         (),                                                                                       // (terminated)
		.in_channel        (1'b0),                                                                                   // (terminated)
		.out_channel       ()                                                                                        // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (77),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (57),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (58),
		.PKT_TRANS_POSTED          (59),
		.PKT_TRANS_WRITE           (60),
		.PKT_TRANS_READ            (61),
		.PKT_TRANS_LOCK            (62),
		.PKT_SRC_ID_H              (85),
		.PKT_SRC_ID_L              (79),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (86),
		.PKT_BURSTWRAP_H           (69),
		.PKT_BURSTWRAP_L           (67),
		.PKT_BYTE_CNT_H            (66),
		.PKT_BYTE_CNT_L            (64),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (72),
		.PKT_BURST_SIZE_L          (70),
		.ST_CHANNEL_W              (99),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) ch3_yn1_u_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                           //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                //       clk_reset.reset
		.m0_address              (ch3_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ch3_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ch3_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ch3_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ch3_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ch3_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ch3_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ch3_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ch3_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ch3_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ch3_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ch3_yn1_u_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ch3_yn1_u_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ch3_yn1_u_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ch3_yn1_u_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ch3_yn1_u_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src69_ready),                                                    //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src69_valid),                                                    //                .valid
		.cp_data                 (cmd_xbar_demux_001_src69_data),                                                     //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src69_startofpacket),                                            //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src69_endofpacket),                                              //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src69_channel),                                                  //                .channel
		.rf_sink_ready           (ch3_yn1_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ch3_yn1_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ch3_yn1_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ch3_yn1_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ch3_yn1_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ch3_yn1_u_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ch3_yn1_u_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ch3_yn1_u_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ch3_yn1_u_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ch3_yn1_u_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ch3_yn1_u_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ch3_yn1_u_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (ch3_yn1_u_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (ch3_yn1_u_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ch3_yn1_u_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ch3_yn1_u_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                             //     (terminated)
		.m0_writeresponserequest (),                                                                                  //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                               //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ch3_yn1_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                           //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                // clk_reset.reset
		.in_data           (ch3_yn1_u_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ch3_yn1_u_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ch3_yn1_u_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ch3_yn1_u_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ch3_yn1_u_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ch3_yn1_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ch3_yn1_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ch3_yn1_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ch3_yn1_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ch3_yn1_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                             // (terminated)
		.csr_read          (1'b0),                                                                              // (terminated)
		.csr_write         (1'b0),                                                                              // (terminated)
		.csr_readdata      (),                                                                                  // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                              // (terminated)
		.almost_full_data  (),                                                                                  // (terminated)
		.almost_empty_data (),                                                                                  // (terminated)
		.in_empty          (1'b0),                                                                              // (terminated)
		.out_empty         (),                                                                                  // (terminated)
		.in_error          (1'b0),                                                                              // (terminated)
		.out_error         (),                                                                                  // (terminated)
		.in_channel        (1'b0),                                                                              // (terminated)
		.out_channel       ()                                                                                   // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (77),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (57),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (58),
		.PKT_TRANS_POSTED          (59),
		.PKT_TRANS_WRITE           (60),
		.PKT_TRANS_READ            (61),
		.PKT_TRANS_LOCK            (62),
		.PKT_SRC_ID_H              (85),
		.PKT_SRC_ID_L              (79),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (86),
		.PKT_BURSTWRAP_H           (69),
		.PKT_BURSTWRAP_L           (67),
		.PKT_BYTE_CNT_H            (66),
		.PKT_BYTE_CNT_L            (64),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (72),
		.PKT_BURST_SIZE_L          (70),
		.ST_CHANNEL_W              (99),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) ch3_time_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                          //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                               //       clk_reset.reset
		.m0_address              (ch3_time_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ch3_time_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ch3_time_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ch3_time_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ch3_time_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ch3_time_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ch3_time_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ch3_time_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ch3_time_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ch3_time_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ch3_time_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ch3_time_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ch3_time_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ch3_time_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ch3_time_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ch3_time_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src70_ready),                                                   //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src70_valid),                                                   //                .valid
		.cp_data                 (cmd_xbar_demux_001_src70_data),                                                    //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src70_startofpacket),                                           //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src70_endofpacket),                                             //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src70_channel),                                                 //                .channel
		.rf_sink_ready           (ch3_time_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ch3_time_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ch3_time_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ch3_time_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ch3_time_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ch3_time_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ch3_time_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ch3_time_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ch3_time_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ch3_time_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ch3_time_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ch3_time_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (ch3_time_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (ch3_time_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ch3_time_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ch3_time_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                            //     (terminated)
		.m0_writeresponserequest (),                                                                                 //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                              //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ch3_time_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                          //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                               // clk_reset.reset
		.in_data           (ch3_time_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ch3_time_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ch3_time_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ch3_time_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ch3_time_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ch3_time_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ch3_time_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ch3_time_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ch3_time_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ch3_time_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                            // (terminated)
		.csr_read          (1'b0),                                                                             // (terminated)
		.csr_write         (1'b0),                                                                             // (terminated)
		.csr_readdata      (),                                                                                 // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                             // (terminated)
		.almost_full_data  (),                                                                                 // (terminated)
		.almost_empty_data (),                                                                                 // (terminated)
		.in_empty          (1'b0),                                                                             // (terminated)
		.out_empty         (),                                                                                 // (terminated)
		.in_error          (1'b0),                                                                             // (terminated)
		.out_error         (),                                                                                 // (terminated)
		.in_channel        (1'b0),                                                                             // (terminated)
		.out_channel       ()                                                                                  // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (77),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (57),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (58),
		.PKT_TRANS_POSTED          (59),
		.PKT_TRANS_WRITE           (60),
		.PKT_TRANS_READ            (61),
		.PKT_TRANS_LOCK            (62),
		.PKT_SRC_ID_H              (85),
		.PKT_SRC_ID_L              (79),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (86),
		.PKT_BURSTWRAP_H           (69),
		.PKT_BURSTWRAP_L           (67),
		.PKT_BYTE_CNT_H            (66),
		.PKT_BYTE_CNT_L            (64),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (72),
		.PKT_BURST_SIZE_L          (70),
		.ST_CHANNEL_W              (99),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) ch3_yn3_l_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                           //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                //       clk_reset.reset
		.m0_address              (ch3_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ch3_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ch3_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ch3_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ch3_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ch3_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ch3_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ch3_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ch3_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ch3_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ch3_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ch3_yn3_l_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ch3_yn3_l_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ch3_yn3_l_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ch3_yn3_l_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ch3_yn3_l_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src71_ready),                                                    //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src71_valid),                                                    //                .valid
		.cp_data                 (cmd_xbar_demux_001_src71_data),                                                     //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src71_startofpacket),                                            //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src71_endofpacket),                                              //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src71_channel),                                                  //                .channel
		.rf_sink_ready           (ch3_yn3_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ch3_yn3_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ch3_yn3_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ch3_yn3_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ch3_yn3_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ch3_yn3_l_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ch3_yn3_l_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ch3_yn3_l_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ch3_yn3_l_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ch3_yn3_l_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ch3_yn3_l_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ch3_yn3_l_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (ch3_yn3_l_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (ch3_yn3_l_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ch3_yn3_l_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ch3_yn3_l_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                             //     (terminated)
		.m0_writeresponserequest (),                                                                                  //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                               //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ch3_yn3_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                           //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                // clk_reset.reset
		.in_data           (ch3_yn3_l_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ch3_yn3_l_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ch3_yn3_l_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ch3_yn3_l_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ch3_yn3_l_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ch3_yn3_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ch3_yn3_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ch3_yn3_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ch3_yn3_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ch3_yn3_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                             // (terminated)
		.csr_read          (1'b0),                                                                              // (terminated)
		.csr_write         (1'b0),                                                                              // (terminated)
		.csr_readdata      (),                                                                                  // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                              // (terminated)
		.almost_full_data  (),                                                                                  // (terminated)
		.almost_empty_data (),                                                                                  // (terminated)
		.in_empty          (1'b0),                                                                              // (terminated)
		.out_empty         (),                                                                                  // (terminated)
		.in_error          (1'b0),                                                                              // (terminated)
		.out_error         (),                                                                                  // (terminated)
		.in_channel        (1'b0),                                                                              // (terminated)
		.out_channel       ()                                                                                   // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (77),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (57),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (58),
		.PKT_TRANS_POSTED          (59),
		.PKT_TRANS_WRITE           (60),
		.PKT_TRANS_READ            (61),
		.PKT_TRANS_LOCK            (62),
		.PKT_SRC_ID_H              (85),
		.PKT_SRC_ID_L              (79),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (86),
		.PKT_BURSTWRAP_H           (69),
		.PKT_BURSTWRAP_L           (67),
		.PKT_BYTE_CNT_H            (66),
		.PKT_BYTE_CNT_L            (64),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (72),
		.PKT_BURST_SIZE_L          (70),
		.ST_CHANNEL_W              (99),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) ch3_yn3_ml_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                            //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                 //       clk_reset.reset
		.m0_address              (ch3_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ch3_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ch3_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ch3_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ch3_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ch3_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ch3_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ch3_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ch3_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ch3_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ch3_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ch3_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ch3_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ch3_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ch3_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ch3_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src72_ready),                                                     //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src72_valid),                                                     //                .valid
		.cp_data                 (cmd_xbar_demux_001_src72_data),                                                      //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src72_startofpacket),                                             //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src72_endofpacket),                                               //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src72_channel),                                                   //                .channel
		.rf_sink_ready           (ch3_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ch3_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ch3_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ch3_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ch3_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ch3_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ch3_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ch3_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ch3_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ch3_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ch3_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ch3_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (ch3_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (ch3_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ch3_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ch3_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                              //     (terminated)
		.m0_writeresponserequest (),                                                                                   //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ch3_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                            //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                 // clk_reset.reset
		.in_data           (ch3_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ch3_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ch3_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ch3_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ch3_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ch3_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ch3_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ch3_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ch3_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ch3_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                              // (terminated)
		.csr_read          (1'b0),                                                                               // (terminated)
		.csr_write         (1'b0),                                                                               // (terminated)
		.csr_readdata      (),                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                               // (terminated)
		.almost_full_data  (),                                                                                   // (terminated)
		.almost_empty_data (),                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                               // (terminated)
		.out_empty         (),                                                                                   // (terminated)
		.in_error          (1'b0),                                                                               // (terminated)
		.out_error         (),                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                               // (terminated)
		.out_channel       ()                                                                                    // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (77),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (57),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (58),
		.PKT_TRANS_POSTED          (59),
		.PKT_TRANS_WRITE           (60),
		.PKT_TRANS_READ            (61),
		.PKT_TRANS_LOCK            (62),
		.PKT_SRC_ID_H              (85),
		.PKT_SRC_ID_L              (79),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (86),
		.PKT_BURSTWRAP_H           (69),
		.PKT_BURSTWRAP_L           (67),
		.PKT_BYTE_CNT_H            (66),
		.PKT_BYTE_CNT_L            (64),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (72),
		.PKT_BURST_SIZE_L          (70),
		.ST_CHANNEL_W              (99),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) ch3_yn3_mu_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                            //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                 //       clk_reset.reset
		.m0_address              (ch3_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ch3_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ch3_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ch3_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ch3_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ch3_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ch3_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ch3_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ch3_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ch3_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ch3_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ch3_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ch3_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ch3_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ch3_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ch3_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src73_ready),                                                     //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src73_valid),                                                     //                .valid
		.cp_data                 (cmd_xbar_demux_001_src73_data),                                                      //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src73_startofpacket),                                             //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src73_endofpacket),                                               //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src73_channel),                                                   //                .channel
		.rf_sink_ready           (ch3_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ch3_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ch3_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ch3_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ch3_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ch3_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ch3_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ch3_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ch3_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ch3_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ch3_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ch3_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (ch3_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (ch3_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ch3_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ch3_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                              //     (terminated)
		.m0_writeresponserequest (),                                                                                   //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ch3_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                            //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                 // clk_reset.reset
		.in_data           (ch3_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ch3_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ch3_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ch3_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ch3_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ch3_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ch3_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ch3_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ch3_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ch3_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                              // (terminated)
		.csr_read          (1'b0),                                                                               // (terminated)
		.csr_write         (1'b0),                                                                               // (terminated)
		.csr_readdata      (),                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                               // (terminated)
		.almost_full_data  (),                                                                                   // (terminated)
		.almost_empty_data (),                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                               // (terminated)
		.out_empty         (),                                                                                   // (terminated)
		.in_error          (1'b0),                                                                               // (terminated)
		.out_error         (),                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                               // (terminated)
		.out_channel       ()                                                                                    // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (77),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (57),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (58),
		.PKT_TRANS_POSTED          (59),
		.PKT_TRANS_WRITE           (60),
		.PKT_TRANS_READ            (61),
		.PKT_TRANS_LOCK            (62),
		.PKT_SRC_ID_H              (85),
		.PKT_SRC_ID_L              (79),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (86),
		.PKT_BURSTWRAP_H           (69),
		.PKT_BURSTWRAP_L           (67),
		.PKT_BYTE_CNT_H            (66),
		.PKT_BYTE_CNT_L            (64),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (72),
		.PKT_BURST_SIZE_L          (70),
		.ST_CHANNEL_W              (99),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) ch3_yn3_u_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                           //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                //       clk_reset.reset
		.m0_address              (ch3_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ch3_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ch3_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ch3_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ch3_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ch3_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ch3_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ch3_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ch3_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ch3_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ch3_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ch3_yn3_u_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ch3_yn3_u_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ch3_yn3_u_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ch3_yn3_u_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ch3_yn3_u_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src74_ready),                                                    //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src74_valid),                                                    //                .valid
		.cp_data                 (cmd_xbar_demux_001_src74_data),                                                     //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src74_startofpacket),                                            //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src74_endofpacket),                                              //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src74_channel),                                                  //                .channel
		.rf_sink_ready           (ch3_yn3_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ch3_yn3_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ch3_yn3_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ch3_yn3_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ch3_yn3_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ch3_yn3_u_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ch3_yn3_u_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ch3_yn3_u_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ch3_yn3_u_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ch3_yn3_u_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ch3_yn3_u_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ch3_yn3_u_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (ch3_yn3_u_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (ch3_yn3_u_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ch3_yn3_u_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ch3_yn3_u_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                             //     (terminated)
		.m0_writeresponserequest (),                                                                                  //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                               //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ch3_yn3_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                           //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                // clk_reset.reset
		.in_data           (ch3_yn3_u_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ch3_yn3_u_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ch3_yn3_u_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ch3_yn3_u_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ch3_yn3_u_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ch3_yn3_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ch3_yn3_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ch3_yn3_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ch3_yn3_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ch3_yn3_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                             // (terminated)
		.csr_read          (1'b0),                                                                              // (terminated)
		.csr_write         (1'b0),                                                                              // (terminated)
		.csr_readdata      (),                                                                                  // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                              // (terminated)
		.almost_full_data  (),                                                                                  // (terminated)
		.almost_empty_data (),                                                                                  // (terminated)
		.in_empty          (1'b0),                                                                              // (terminated)
		.out_empty         (),                                                                                  // (terminated)
		.in_error          (1'b0),                                                                              // (terminated)
		.out_error         (),                                                                                  // (terminated)
		.in_channel        (1'b0),                                                                              // (terminated)
		.out_channel       ()                                                                                   // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (77),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (57),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (58),
		.PKT_TRANS_POSTED          (59),
		.PKT_TRANS_WRITE           (60),
		.PKT_TRANS_READ            (61),
		.PKT_TRANS_LOCK            (62),
		.PKT_SRC_ID_H              (85),
		.PKT_SRC_ID_L              (79),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (86),
		.PKT_BURSTWRAP_H           (69),
		.PKT_BURSTWRAP_L           (67),
		.PKT_BYTE_CNT_H            (66),
		.PKT_BYTE_CNT_L            (64),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (72),
		.PKT_BURST_SIZE_L          (70),
		.ST_CHANNEL_W              (99),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) ch3_yn2_l_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                           //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                //       clk_reset.reset
		.m0_address              (ch3_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ch3_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ch3_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ch3_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ch3_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ch3_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ch3_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ch3_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ch3_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ch3_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ch3_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ch3_yn2_l_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ch3_yn2_l_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ch3_yn2_l_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ch3_yn2_l_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ch3_yn2_l_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src75_ready),                                                    //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src75_valid),                                                    //                .valid
		.cp_data                 (cmd_xbar_demux_001_src75_data),                                                     //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src75_startofpacket),                                            //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src75_endofpacket),                                              //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src75_channel),                                                  //                .channel
		.rf_sink_ready           (ch3_yn2_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ch3_yn2_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ch3_yn2_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ch3_yn2_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ch3_yn2_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ch3_yn2_l_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ch3_yn2_l_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ch3_yn2_l_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ch3_yn2_l_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ch3_yn2_l_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ch3_yn2_l_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ch3_yn2_l_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (ch3_yn2_l_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (ch3_yn2_l_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ch3_yn2_l_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ch3_yn2_l_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                             //     (terminated)
		.m0_writeresponserequest (),                                                                                  //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                               //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ch3_yn2_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                           //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                // clk_reset.reset
		.in_data           (ch3_yn2_l_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ch3_yn2_l_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ch3_yn2_l_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ch3_yn2_l_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ch3_yn2_l_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ch3_yn2_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ch3_yn2_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ch3_yn2_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ch3_yn2_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ch3_yn2_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                             // (terminated)
		.csr_read          (1'b0),                                                                              // (terminated)
		.csr_write         (1'b0),                                                                              // (terminated)
		.csr_readdata      (),                                                                                  // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                              // (terminated)
		.almost_full_data  (),                                                                                  // (terminated)
		.almost_empty_data (),                                                                                  // (terminated)
		.in_empty          (1'b0),                                                                              // (terminated)
		.out_empty         (),                                                                                  // (terminated)
		.in_error          (1'b0),                                                                              // (terminated)
		.out_error         (),                                                                                  // (terminated)
		.in_channel        (1'b0),                                                                              // (terminated)
		.out_channel       ()                                                                                   // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (77),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (57),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (58),
		.PKT_TRANS_POSTED          (59),
		.PKT_TRANS_WRITE           (60),
		.PKT_TRANS_READ            (61),
		.PKT_TRANS_LOCK            (62),
		.PKT_SRC_ID_H              (85),
		.PKT_SRC_ID_L              (79),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (86),
		.PKT_BURSTWRAP_H           (69),
		.PKT_BURSTWRAP_L           (67),
		.PKT_BYTE_CNT_H            (66),
		.PKT_BYTE_CNT_L            (64),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (72),
		.PKT_BURST_SIZE_L          (70),
		.ST_CHANNEL_W              (99),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) ch3_yn2_ml_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                            //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                 //       clk_reset.reset
		.m0_address              (ch3_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ch3_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ch3_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ch3_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ch3_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ch3_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ch3_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ch3_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ch3_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ch3_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ch3_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ch3_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ch3_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ch3_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ch3_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ch3_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src76_ready),                                                     //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src76_valid),                                                     //                .valid
		.cp_data                 (cmd_xbar_demux_001_src76_data),                                                      //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src76_startofpacket),                                             //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src76_endofpacket),                                               //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src76_channel),                                                   //                .channel
		.rf_sink_ready           (ch3_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ch3_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ch3_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ch3_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ch3_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ch3_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ch3_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ch3_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ch3_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ch3_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ch3_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ch3_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (ch3_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (ch3_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ch3_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ch3_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                              //     (terminated)
		.m0_writeresponserequest (),                                                                                   //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ch3_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                            //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                 // clk_reset.reset
		.in_data           (ch3_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ch3_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ch3_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ch3_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ch3_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ch3_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ch3_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ch3_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ch3_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ch3_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                              // (terminated)
		.csr_read          (1'b0),                                                                               // (terminated)
		.csr_write         (1'b0),                                                                               // (terminated)
		.csr_readdata      (),                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                               // (terminated)
		.almost_full_data  (),                                                                                   // (terminated)
		.almost_empty_data (),                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                               // (terminated)
		.out_empty         (),                                                                                   // (terminated)
		.in_error          (1'b0),                                                                               // (terminated)
		.out_error         (),                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                               // (terminated)
		.out_channel       ()                                                                                    // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (77),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (57),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (58),
		.PKT_TRANS_POSTED          (59),
		.PKT_TRANS_WRITE           (60),
		.PKT_TRANS_READ            (61),
		.PKT_TRANS_LOCK            (62),
		.PKT_SRC_ID_H              (85),
		.PKT_SRC_ID_L              (79),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (86),
		.PKT_BURSTWRAP_H           (69),
		.PKT_BURSTWRAP_L           (67),
		.PKT_BYTE_CNT_H            (66),
		.PKT_BYTE_CNT_L            (64),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (72),
		.PKT_BURST_SIZE_L          (70),
		.ST_CHANNEL_W              (99),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) ch3_yn2_mu_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                            //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                 //       clk_reset.reset
		.m0_address              (ch3_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ch3_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ch3_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ch3_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ch3_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ch3_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ch3_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ch3_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ch3_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ch3_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ch3_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ch3_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ch3_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ch3_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ch3_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ch3_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src77_ready),                                                     //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src77_valid),                                                     //                .valid
		.cp_data                 (cmd_xbar_demux_001_src77_data),                                                      //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src77_startofpacket),                                             //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src77_endofpacket),                                               //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src77_channel),                                                   //                .channel
		.rf_sink_ready           (ch3_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ch3_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ch3_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ch3_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ch3_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ch3_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ch3_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ch3_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ch3_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ch3_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ch3_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ch3_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (ch3_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (ch3_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ch3_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ch3_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                              //     (terminated)
		.m0_writeresponserequest (),                                                                                   //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ch3_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                            //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                 // clk_reset.reset
		.in_data           (ch3_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ch3_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ch3_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ch3_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ch3_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ch3_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ch3_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ch3_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ch3_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ch3_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                              // (terminated)
		.csr_read          (1'b0),                                                                               // (terminated)
		.csr_write         (1'b0),                                                                               // (terminated)
		.csr_readdata      (),                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                               // (terminated)
		.almost_full_data  (),                                                                                   // (terminated)
		.almost_empty_data (),                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                               // (terminated)
		.out_empty         (),                                                                                   // (terminated)
		.in_error          (1'b0),                                                                               // (terminated)
		.out_error         (),                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                               // (terminated)
		.out_channel       ()                                                                                    // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (77),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (57),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (58),
		.PKT_TRANS_POSTED          (59),
		.PKT_TRANS_WRITE           (60),
		.PKT_TRANS_READ            (61),
		.PKT_TRANS_LOCK            (62),
		.PKT_SRC_ID_H              (85),
		.PKT_SRC_ID_L              (79),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (86),
		.PKT_BURSTWRAP_H           (69),
		.PKT_BURSTWRAP_L           (67),
		.PKT_BYTE_CNT_H            (66),
		.PKT_BYTE_CNT_L            (64),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (72),
		.PKT_BURST_SIZE_L          (70),
		.ST_CHANNEL_W              (99),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) ch3_yn2_u_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                           //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                //       clk_reset.reset
		.m0_address              (ch3_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ch3_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ch3_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ch3_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ch3_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ch3_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ch3_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ch3_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ch3_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ch3_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ch3_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ch3_yn2_u_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ch3_yn2_u_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ch3_yn2_u_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ch3_yn2_u_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ch3_yn2_u_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src78_ready),                                                    //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src78_valid),                                                    //                .valid
		.cp_data                 (cmd_xbar_demux_001_src78_data),                                                     //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src78_startofpacket),                                            //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src78_endofpacket),                                              //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src78_channel),                                                  //                .channel
		.rf_sink_ready           (ch3_yn2_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ch3_yn2_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ch3_yn2_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ch3_yn2_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ch3_yn2_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ch3_yn2_u_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ch3_yn2_u_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ch3_yn2_u_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ch3_yn2_u_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ch3_yn2_u_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ch3_yn2_u_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ch3_yn2_u_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (ch3_yn2_u_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (ch3_yn2_u_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ch3_yn2_u_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ch3_yn2_u_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                             //     (terminated)
		.m0_writeresponserequest (),                                                                                  //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                               //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ch3_yn2_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                           //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                // clk_reset.reset
		.in_data           (ch3_yn2_u_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ch3_yn2_u_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ch3_yn2_u_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ch3_yn2_u_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ch3_yn2_u_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ch3_yn2_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ch3_yn2_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ch3_yn2_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ch3_yn2_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ch3_yn2_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                             // (terminated)
		.csr_read          (1'b0),                                                                              // (terminated)
		.csr_write         (1'b0),                                                                              // (terminated)
		.csr_readdata      (),                                                                                  // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                              // (terminated)
		.almost_full_data  (),                                                                                  // (terminated)
		.almost_empty_data (),                                                                                  // (terminated)
		.in_empty          (1'b0),                                                                              // (terminated)
		.out_empty         (),                                                                                  // (terminated)
		.in_error          (1'b0),                                                                              // (terminated)
		.out_error         (),                                                                                  // (terminated)
		.in_channel        (1'b0),                                                                              // (terminated)
		.out_channel       ()                                                                                   // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (77),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (57),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (58),
		.PKT_TRANS_POSTED          (59),
		.PKT_TRANS_WRITE           (60),
		.PKT_TRANS_READ            (61),
		.PKT_TRANS_LOCK            (62),
		.PKT_SRC_ID_H              (85),
		.PKT_SRC_ID_L              (79),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (86),
		.PKT_BURSTWRAP_H           (69),
		.PKT_BURSTWRAP_L           (67),
		.PKT_BYTE_CNT_H            (66),
		.PKT_BYTE_CNT_L            (64),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (72),
		.PKT_BURST_SIZE_L          (70),
		.ST_CHANNEL_W              (99),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) ch3_yn1_l_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                           //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                //       clk_reset.reset
		.m0_address              (ch3_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ch3_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ch3_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ch3_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ch3_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ch3_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ch3_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ch3_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ch3_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ch3_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ch3_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ch3_yn1_l_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ch3_yn1_l_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ch3_yn1_l_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ch3_yn1_l_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ch3_yn1_l_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src79_ready),                                                    //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src79_valid),                                                    //                .valid
		.cp_data                 (cmd_xbar_demux_001_src79_data),                                                     //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src79_startofpacket),                                            //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src79_endofpacket),                                              //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src79_channel),                                                  //                .channel
		.rf_sink_ready           (ch3_yn1_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ch3_yn1_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ch3_yn1_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ch3_yn1_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ch3_yn1_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ch3_yn1_l_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ch3_yn1_l_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ch3_yn1_l_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ch3_yn1_l_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ch3_yn1_l_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ch3_yn1_l_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ch3_yn1_l_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (ch3_yn1_l_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (ch3_yn1_l_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ch3_yn1_l_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ch3_yn1_l_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                             //     (terminated)
		.m0_writeresponserequest (),                                                                                  //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                               //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ch3_yn1_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                           //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                // clk_reset.reset
		.in_data           (ch3_yn1_l_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ch3_yn1_l_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ch3_yn1_l_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ch3_yn1_l_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ch3_yn1_l_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ch3_yn1_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ch3_yn1_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ch3_yn1_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ch3_yn1_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ch3_yn1_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                             // (terminated)
		.csr_read          (1'b0),                                                                              // (terminated)
		.csr_write         (1'b0),                                                                              // (terminated)
		.csr_readdata      (),                                                                                  // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                              // (terminated)
		.almost_full_data  (),                                                                                  // (terminated)
		.almost_empty_data (),                                                                                  // (terminated)
		.in_empty          (1'b0),                                                                              // (terminated)
		.out_empty         (),                                                                                  // (terminated)
		.in_error          (1'b0),                                                                              // (terminated)
		.out_error         (),                                                                                  // (terminated)
		.in_channel        (1'b0),                                                                              // (terminated)
		.out_channel       ()                                                                                   // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (77),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (57),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (58),
		.PKT_TRANS_POSTED          (59),
		.PKT_TRANS_WRITE           (60),
		.PKT_TRANS_READ            (61),
		.PKT_TRANS_LOCK            (62),
		.PKT_SRC_ID_H              (85),
		.PKT_SRC_ID_L              (79),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (86),
		.PKT_BURSTWRAP_H           (69),
		.PKT_BURSTWRAP_L           (67),
		.PKT_BYTE_CNT_H            (66),
		.PKT_BYTE_CNT_L            (64),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (72),
		.PKT_BURST_SIZE_L          (70),
		.ST_CHANNEL_W              (99),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) ch3_yn1_mu_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                            //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                 //       clk_reset.reset
		.m0_address              (ch3_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ch3_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ch3_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ch3_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ch3_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ch3_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ch3_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ch3_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ch3_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ch3_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ch3_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ch3_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ch3_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ch3_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ch3_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ch3_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src80_ready),                                                     //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src80_valid),                                                     //                .valid
		.cp_data                 (cmd_xbar_demux_001_src80_data),                                                      //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src80_startofpacket),                                             //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src80_endofpacket),                                               //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src80_channel),                                                   //                .channel
		.rf_sink_ready           (ch3_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ch3_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ch3_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ch3_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ch3_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ch3_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ch3_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ch3_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ch3_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ch3_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ch3_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ch3_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (ch3_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (ch3_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ch3_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ch3_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                              //     (terminated)
		.m0_writeresponserequest (),                                                                                   //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ch3_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                            //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                 // clk_reset.reset
		.in_data           (ch3_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ch3_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ch3_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ch3_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ch3_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ch3_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ch3_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ch3_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ch3_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ch3_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                              // (terminated)
		.csr_read          (1'b0),                                                                               // (terminated)
		.csr_write         (1'b0),                                                                               // (terminated)
		.csr_readdata      (),                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                               // (terminated)
		.almost_full_data  (),                                                                                   // (terminated)
		.almost_empty_data (),                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                               // (terminated)
		.out_empty         (),                                                                                   // (terminated)
		.in_error          (1'b0),                                                                               // (terminated)
		.out_error         (),                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                               // (terminated)
		.out_channel       ()                                                                                    // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (77),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (57),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (58),
		.PKT_TRANS_POSTED          (59),
		.PKT_TRANS_WRITE           (60),
		.PKT_TRANS_READ            (61),
		.PKT_TRANS_LOCK            (62),
		.PKT_SRC_ID_H              (85),
		.PKT_SRC_ID_L              (79),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (86),
		.PKT_BURSTWRAP_H           (69),
		.PKT_BURSTWRAP_L           (67),
		.PKT_BYTE_CNT_H            (66),
		.PKT_BYTE_CNT_L            (64),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (72),
		.PKT_BURST_SIZE_L          (70),
		.ST_CHANNEL_W              (99),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) ch3_yn1_ml_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                            //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                 //       clk_reset.reset
		.m0_address              (ch3_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ch3_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ch3_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ch3_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ch3_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ch3_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ch3_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ch3_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ch3_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ch3_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ch3_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ch3_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ch3_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ch3_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ch3_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ch3_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src81_ready),                                                     //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src81_valid),                                                     //                .valid
		.cp_data                 (cmd_xbar_demux_001_src81_data),                                                      //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src81_startofpacket),                                             //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src81_endofpacket),                                               //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src81_channel),                                                   //                .channel
		.rf_sink_ready           (ch3_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ch3_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ch3_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ch3_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ch3_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ch3_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ch3_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ch3_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ch3_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ch3_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ch3_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ch3_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (ch3_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (ch3_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ch3_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ch3_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                              //     (terminated)
		.m0_writeresponserequest (),                                                                                   //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ch3_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                            //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                 // clk_reset.reset
		.in_data           (ch3_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ch3_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ch3_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ch3_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ch3_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ch3_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ch3_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ch3_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ch3_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ch3_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                              // (terminated)
		.csr_read          (1'b0),                                                                               // (terminated)
		.csr_write         (1'b0),                                                                               // (terminated)
		.csr_readdata      (),                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                               // (terminated)
		.almost_full_data  (),                                                                                   // (terminated)
		.almost_empty_data (),                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                               // (terminated)
		.out_empty         (),                                                                                   // (terminated)
		.in_error          (1'b0),                                                                               // (terminated)
		.out_error         (),                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                               // (terminated)
		.out_channel       ()                                                                                    // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (77),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (57),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (58),
		.PKT_TRANS_POSTED          (59),
		.PKT_TRANS_WRITE           (60),
		.PKT_TRANS_READ            (61),
		.PKT_TRANS_LOCK            (62),
		.PKT_SRC_ID_H              (85),
		.PKT_SRC_ID_L              (79),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (86),
		.PKT_BURSTWRAP_H           (69),
		.PKT_BURSTWRAP_L           (67),
		.PKT_BYTE_CNT_H            (66),
		.PKT_BYTE_CNT_L            (64),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (72),
		.PKT_BURST_SIZE_L          (70),
		.ST_CHANNEL_W              (99),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) ch4_timer_rst_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                               //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                    //       clk_reset.reset
		.m0_address              (ch4_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ch4_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ch4_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ch4_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ch4_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ch4_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ch4_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ch4_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ch4_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ch4_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ch4_timer_rst_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ch4_timer_rst_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ch4_timer_rst_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ch4_timer_rst_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ch4_timer_rst_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ch4_timer_rst_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src82_ready),                                                        //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src82_valid),                                                        //                .valid
		.cp_data                 (cmd_xbar_demux_001_src82_data),                                                         //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src82_startofpacket),                                                //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src82_endofpacket),                                                  //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src82_channel),                                                      //                .channel
		.rf_sink_ready           (ch4_timer_rst_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ch4_timer_rst_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ch4_timer_rst_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ch4_timer_rst_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ch4_timer_rst_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ch4_timer_rst_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ch4_timer_rst_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ch4_timer_rst_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ch4_timer_rst_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ch4_timer_rst_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ch4_timer_rst_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ch4_timer_rst_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (ch4_timer_rst_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (ch4_timer_rst_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ch4_timer_rst_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ch4_timer_rst_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                 //     (terminated)
		.m0_writeresponserequest (),                                                                                      //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                   //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ch4_timer_rst_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                               //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                    // clk_reset.reset
		.in_data           (ch4_timer_rst_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ch4_timer_rst_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ch4_timer_rst_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ch4_timer_rst_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ch4_timer_rst_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ch4_timer_rst_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ch4_timer_rst_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ch4_timer_rst_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ch4_timer_rst_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ch4_timer_rst_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                 // (terminated)
		.csr_read          (1'b0),                                                                                  // (terminated)
		.csr_write         (1'b0),                                                                                  // (terminated)
		.csr_readdata      (),                                                                                      // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                  // (terminated)
		.almost_full_data  (),                                                                                      // (terminated)
		.almost_empty_data (),                                                                                      // (terminated)
		.in_empty          (1'b0),                                                                                  // (terminated)
		.out_empty         (),                                                                                      // (terminated)
		.in_error          (1'b0),                                                                                  // (terminated)
		.out_error         (),                                                                                      // (terminated)
		.in_channel        (1'b0),                                                                                  // (terminated)
		.out_channel       ()                                                                                       // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (77),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (57),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (58),
		.PKT_TRANS_POSTED          (59),
		.PKT_TRANS_WRITE           (60),
		.PKT_TRANS_READ            (61),
		.PKT_TRANS_LOCK            (62),
		.PKT_SRC_ID_H              (85),
		.PKT_SRC_ID_L              (79),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (86),
		.PKT_BURSTWRAP_H           (69),
		.PKT_BURSTWRAP_L           (67),
		.PKT_BYTE_CNT_H            (66),
		.PKT_BYTE_CNT_L            (64),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (72),
		.PKT_BURST_SIZE_L          (70),
		.ST_CHANNEL_W              (99),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) ch4_thresh_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                            //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                 //       clk_reset.reset
		.m0_address              (ch4_thresh_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ch4_thresh_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ch4_thresh_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ch4_thresh_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ch4_thresh_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ch4_thresh_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ch4_thresh_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ch4_thresh_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ch4_thresh_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ch4_thresh_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ch4_thresh_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ch4_thresh_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ch4_thresh_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ch4_thresh_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ch4_thresh_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ch4_thresh_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src83_ready),                                                     //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src83_valid),                                                     //                .valid
		.cp_data                 (cmd_xbar_demux_001_src83_data),                                                      //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src83_startofpacket),                                             //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src83_endofpacket),                                               //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src83_channel),                                                   //                .channel
		.rf_sink_ready           (ch4_thresh_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ch4_thresh_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ch4_thresh_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ch4_thresh_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ch4_thresh_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ch4_thresh_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ch4_thresh_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ch4_thresh_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ch4_thresh_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ch4_thresh_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ch4_thresh_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ch4_thresh_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (ch4_thresh_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (ch4_thresh_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ch4_thresh_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ch4_thresh_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                              //     (terminated)
		.m0_writeresponserequest (),                                                                                   //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ch4_thresh_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                            //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                 // clk_reset.reset
		.in_data           (ch4_thresh_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ch4_thresh_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ch4_thresh_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ch4_thresh_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ch4_thresh_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ch4_thresh_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ch4_thresh_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ch4_thresh_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ch4_thresh_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ch4_thresh_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                              // (terminated)
		.csr_read          (1'b0),                                                                               // (terminated)
		.csr_write         (1'b0),                                                                               // (terminated)
		.csr_readdata      (),                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                               // (terminated)
		.almost_full_data  (),                                                                                   // (terminated)
		.almost_empty_data (),                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                               // (terminated)
		.out_empty         (),                                                                                   // (terminated)
		.in_error          (1'b0),                                                                               // (terminated)
		.out_error         (),                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                               // (terminated)
		.out_channel       ()                                                                                    // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (77),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (57),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (58),
		.PKT_TRANS_POSTED          (59),
		.PKT_TRANS_WRITE           (60),
		.PKT_TRANS_READ            (61),
		.PKT_TRANS_LOCK            (62),
		.PKT_SRC_ID_H              (85),
		.PKT_SRC_ID_L              (79),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (86),
		.PKT_BURSTWRAP_H           (69),
		.PKT_BURSTWRAP_L           (67),
		.PKT_BYTE_CNT_H            (66),
		.PKT_BYTE_CNT_L            (64),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (72),
		.PKT_BURST_SIZE_L          (70),
		.ST_CHANNEL_W              (99),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) ch4_rd_peak_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                             //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                  //       clk_reset.reset
		.m0_address              (ch4_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ch4_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ch4_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ch4_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ch4_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ch4_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ch4_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ch4_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ch4_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ch4_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ch4_rd_peak_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ch4_rd_peak_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ch4_rd_peak_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ch4_rd_peak_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ch4_rd_peak_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ch4_rd_peak_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src84_ready),                                                      //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src84_valid),                                                      //                .valid
		.cp_data                 (cmd_xbar_demux_001_src84_data),                                                       //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src84_startofpacket),                                              //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src84_endofpacket),                                                //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src84_channel),                                                    //                .channel
		.rf_sink_ready           (ch4_rd_peak_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ch4_rd_peak_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ch4_rd_peak_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ch4_rd_peak_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ch4_rd_peak_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ch4_rd_peak_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ch4_rd_peak_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ch4_rd_peak_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ch4_rd_peak_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ch4_rd_peak_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ch4_rd_peak_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ch4_rd_peak_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (ch4_rd_peak_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (ch4_rd_peak_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ch4_rd_peak_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ch4_rd_peak_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                               //     (terminated)
		.m0_writeresponserequest (),                                                                                    //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                 //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ch4_rd_peak_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                             //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                  // clk_reset.reset
		.in_data           (ch4_rd_peak_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ch4_rd_peak_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ch4_rd_peak_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ch4_rd_peak_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ch4_rd_peak_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ch4_rd_peak_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ch4_rd_peak_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ch4_rd_peak_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ch4_rd_peak_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ch4_rd_peak_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                               // (terminated)
		.csr_read          (1'b0),                                                                                // (terminated)
		.csr_write         (1'b0),                                                                                // (terminated)
		.csr_readdata      (),                                                                                    // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                // (terminated)
		.almost_full_data  (),                                                                                    // (terminated)
		.almost_empty_data (),                                                                                    // (terminated)
		.in_empty          (1'b0),                                                                                // (terminated)
		.out_empty         (),                                                                                    // (terminated)
		.in_error          (1'b0),                                                                                // (terminated)
		.out_error         (),                                                                                    // (terminated)
		.in_channel        (1'b0),                                                                                // (terminated)
		.out_channel       ()                                                                                     // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (77),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (57),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (58),
		.PKT_TRANS_POSTED          (59),
		.PKT_TRANS_WRITE           (60),
		.PKT_TRANS_READ            (61),
		.PKT_TRANS_LOCK            (62),
		.PKT_SRC_ID_H              (85),
		.PKT_SRC_ID_L              (79),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (86),
		.PKT_BURSTWRAP_H           (69),
		.PKT_BURSTWRAP_L           (67),
		.PKT_BYTE_CNT_H            (66),
		.PKT_BYTE_CNT_L            (64),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (72),
		.PKT_BURST_SIZE_L          (70),
		.ST_CHANNEL_W              (99),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) ch4_peak_found_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                     //       clk_reset.reset
		.m0_address              (ch4_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ch4_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ch4_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ch4_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ch4_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ch4_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ch4_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ch4_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ch4_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ch4_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ch4_peak_found_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ch4_peak_found_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ch4_peak_found_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ch4_peak_found_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ch4_peak_found_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ch4_peak_found_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src85_ready),                                                         //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src85_valid),                                                         //                .valid
		.cp_data                 (cmd_xbar_demux_001_src85_data),                                                          //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src85_startofpacket),                                                 //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src85_endofpacket),                                                   //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src85_channel),                                                       //                .channel
		.rf_sink_ready           (ch4_peak_found_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ch4_peak_found_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ch4_peak_found_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ch4_peak_found_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ch4_peak_found_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ch4_peak_found_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ch4_peak_found_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ch4_peak_found_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ch4_peak_found_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ch4_peak_found_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ch4_peak_found_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ch4_peak_found_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (ch4_peak_found_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (ch4_peak_found_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ch4_peak_found_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ch4_peak_found_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                  //     (terminated)
		.m0_writeresponserequest (),                                                                                       //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                    //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ch4_peak_found_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                     // clk_reset.reset
		.in_data           (ch4_peak_found_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ch4_peak_found_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ch4_peak_found_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ch4_peak_found_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ch4_peak_found_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ch4_peak_found_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ch4_peak_found_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ch4_peak_found_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ch4_peak_found_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ch4_peak_found_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                  // (terminated)
		.csr_read          (1'b0),                                                                                   // (terminated)
		.csr_write         (1'b0),                                                                                   // (terminated)
		.csr_readdata      (),                                                                                       // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                   // (terminated)
		.almost_full_data  (),                                                                                       // (terminated)
		.almost_empty_data (),                                                                                       // (terminated)
		.in_empty          (1'b0),                                                                                   // (terminated)
		.out_empty         (),                                                                                       // (terminated)
		.in_error          (1'b0),                                                                                   // (terminated)
		.out_error         (),                                                                                       // (terminated)
		.in_channel        (1'b0),                                                                                   // (terminated)
		.out_channel       ()                                                                                        // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (77),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (57),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (58),
		.PKT_TRANS_POSTED          (59),
		.PKT_TRANS_WRITE           (60),
		.PKT_TRANS_READ            (61),
		.PKT_TRANS_LOCK            (62),
		.PKT_SRC_ID_H              (85),
		.PKT_SRC_ID_L              (79),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (86),
		.PKT_BURSTWRAP_H           (69),
		.PKT_BURSTWRAP_L           (67),
		.PKT_BYTE_CNT_H            (66),
		.PKT_BYTE_CNT_L            (64),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (72),
		.PKT_BURST_SIZE_L          (70),
		.ST_CHANNEL_W              (99),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) ch4_time_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                          //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                               //       clk_reset.reset
		.m0_address              (ch4_time_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ch4_time_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ch4_time_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ch4_time_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ch4_time_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ch4_time_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ch4_time_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ch4_time_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ch4_time_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ch4_time_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ch4_time_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ch4_time_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ch4_time_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ch4_time_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ch4_time_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ch4_time_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src86_ready),                                                   //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src86_valid),                                                   //                .valid
		.cp_data                 (cmd_xbar_demux_001_src86_data),                                                    //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src86_startofpacket),                                           //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src86_endofpacket),                                             //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src86_channel),                                                 //                .channel
		.rf_sink_ready           (ch4_time_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ch4_time_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ch4_time_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ch4_time_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ch4_time_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ch4_time_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ch4_time_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ch4_time_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ch4_time_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ch4_time_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ch4_time_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ch4_time_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (ch4_time_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (ch4_time_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ch4_time_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ch4_time_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                            //     (terminated)
		.m0_writeresponserequest (),                                                                                 //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                              //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ch4_time_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                          //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                               // clk_reset.reset
		.in_data           (ch4_time_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ch4_time_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ch4_time_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ch4_time_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ch4_time_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ch4_time_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ch4_time_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ch4_time_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ch4_time_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ch4_time_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                            // (terminated)
		.csr_read          (1'b0),                                                                             // (terminated)
		.csr_write         (1'b0),                                                                             // (terminated)
		.csr_readdata      (),                                                                                 // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                             // (terminated)
		.almost_full_data  (),                                                                                 // (terminated)
		.almost_empty_data (),                                                                                 // (terminated)
		.in_empty          (1'b0),                                                                             // (terminated)
		.out_empty         (),                                                                                 // (terminated)
		.in_error          (1'b0),                                                                             // (terminated)
		.out_error         (),                                                                                 // (terminated)
		.in_channel        (1'b0),                                                                             // (terminated)
		.out_channel       ()                                                                                  // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (77),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (57),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (58),
		.PKT_TRANS_POSTED          (59),
		.PKT_TRANS_WRITE           (60),
		.PKT_TRANS_READ            (61),
		.PKT_TRANS_LOCK            (62),
		.PKT_SRC_ID_H              (85),
		.PKT_SRC_ID_L              (79),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (86),
		.PKT_BURSTWRAP_H           (69),
		.PKT_BURSTWRAP_L           (67),
		.PKT_BYTE_CNT_H            (66),
		.PKT_BYTE_CNT_L            (64),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (72),
		.PKT_BURST_SIZE_L          (70),
		.ST_CHANNEL_W              (99),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) ch4_yn1_u_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                           //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                //       clk_reset.reset
		.m0_address              (ch4_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ch4_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ch4_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ch4_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ch4_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ch4_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ch4_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ch4_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ch4_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ch4_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ch4_yn1_u_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ch4_yn1_u_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ch4_yn1_u_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ch4_yn1_u_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ch4_yn1_u_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ch4_yn1_u_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src87_ready),                                                    //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src87_valid),                                                    //                .valid
		.cp_data                 (cmd_xbar_demux_001_src87_data),                                                     //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src87_startofpacket),                                            //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src87_endofpacket),                                              //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src87_channel),                                                  //                .channel
		.rf_sink_ready           (ch4_yn1_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ch4_yn1_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ch4_yn1_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ch4_yn1_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ch4_yn1_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ch4_yn1_u_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ch4_yn1_u_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ch4_yn1_u_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ch4_yn1_u_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ch4_yn1_u_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ch4_yn1_u_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ch4_yn1_u_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (ch4_yn1_u_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (ch4_yn1_u_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ch4_yn1_u_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ch4_yn1_u_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                             //     (terminated)
		.m0_writeresponserequest (),                                                                                  //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                               //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ch4_yn1_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                           //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                // clk_reset.reset
		.in_data           (ch4_yn1_u_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ch4_yn1_u_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ch4_yn1_u_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ch4_yn1_u_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ch4_yn1_u_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ch4_yn1_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ch4_yn1_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ch4_yn1_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ch4_yn1_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ch4_yn1_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                             // (terminated)
		.csr_read          (1'b0),                                                                              // (terminated)
		.csr_write         (1'b0),                                                                              // (terminated)
		.csr_readdata      (),                                                                                  // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                              // (terminated)
		.almost_full_data  (),                                                                                  // (terminated)
		.almost_empty_data (),                                                                                  // (terminated)
		.in_empty          (1'b0),                                                                              // (terminated)
		.out_empty         (),                                                                                  // (terminated)
		.in_error          (1'b0),                                                                              // (terminated)
		.out_error         (),                                                                                  // (terminated)
		.in_channel        (1'b0),                                                                              // (terminated)
		.out_channel       ()                                                                                   // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (77),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (57),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (58),
		.PKT_TRANS_POSTED          (59),
		.PKT_TRANS_WRITE           (60),
		.PKT_TRANS_READ            (61),
		.PKT_TRANS_LOCK            (62),
		.PKT_SRC_ID_H              (85),
		.PKT_SRC_ID_L              (79),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (86),
		.PKT_BURSTWRAP_H           (69),
		.PKT_BURSTWRAP_L           (67),
		.PKT_BYTE_CNT_H            (66),
		.PKT_BYTE_CNT_L            (64),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (72),
		.PKT_BURST_SIZE_L          (70),
		.ST_CHANNEL_W              (99),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) ch4_yn1_mu_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                            //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                 //       clk_reset.reset
		.m0_address              (ch4_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ch4_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ch4_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ch4_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ch4_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ch4_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ch4_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ch4_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ch4_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ch4_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ch4_yn1_mu_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ch4_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ch4_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ch4_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ch4_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ch4_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src88_ready),                                                     //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src88_valid),                                                     //                .valid
		.cp_data                 (cmd_xbar_demux_001_src88_data),                                                      //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src88_startofpacket),                                             //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src88_endofpacket),                                               //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src88_channel),                                                   //                .channel
		.rf_sink_ready           (ch4_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ch4_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ch4_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ch4_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ch4_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ch4_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ch4_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ch4_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ch4_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ch4_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ch4_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ch4_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (ch4_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (ch4_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ch4_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ch4_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                              //     (terminated)
		.m0_writeresponserequest (),                                                                                   //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ch4_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                            //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                 // clk_reset.reset
		.in_data           (ch4_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ch4_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ch4_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ch4_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ch4_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ch4_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ch4_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ch4_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ch4_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ch4_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                              // (terminated)
		.csr_read          (1'b0),                                                                               // (terminated)
		.csr_write         (1'b0),                                                                               // (terminated)
		.csr_readdata      (),                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                               // (terminated)
		.almost_full_data  (),                                                                                   // (terminated)
		.almost_empty_data (),                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                               // (terminated)
		.out_empty         (),                                                                                   // (terminated)
		.in_error          (1'b0),                                                                               // (terminated)
		.out_error         (),                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                               // (terminated)
		.out_channel       ()                                                                                    // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (77),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (57),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (58),
		.PKT_TRANS_POSTED          (59),
		.PKT_TRANS_WRITE           (60),
		.PKT_TRANS_READ            (61),
		.PKT_TRANS_LOCK            (62),
		.PKT_SRC_ID_H              (85),
		.PKT_SRC_ID_L              (79),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (86),
		.PKT_BURSTWRAP_H           (69),
		.PKT_BURSTWRAP_L           (67),
		.PKT_BYTE_CNT_H            (66),
		.PKT_BYTE_CNT_L            (64),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (72),
		.PKT_BURST_SIZE_L          (70),
		.ST_CHANNEL_W              (99),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) ch4_yn1_ml_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                            //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                 //       clk_reset.reset
		.m0_address              (ch4_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ch4_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ch4_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ch4_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ch4_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ch4_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ch4_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ch4_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ch4_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ch4_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ch4_yn1_ml_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ch4_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ch4_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ch4_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ch4_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ch4_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src89_ready),                                                     //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src89_valid),                                                     //                .valid
		.cp_data                 (cmd_xbar_demux_001_src89_data),                                                      //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src89_startofpacket),                                             //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src89_endofpacket),                                               //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src89_channel),                                                   //                .channel
		.rf_sink_ready           (ch4_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ch4_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ch4_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ch4_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ch4_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ch4_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ch4_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ch4_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ch4_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ch4_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ch4_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ch4_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (ch4_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (ch4_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ch4_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ch4_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                              //     (terminated)
		.m0_writeresponserequest (),                                                                                   //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ch4_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                            //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                 // clk_reset.reset
		.in_data           (ch4_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ch4_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ch4_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ch4_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ch4_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ch4_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ch4_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ch4_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ch4_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ch4_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                              // (terminated)
		.csr_read          (1'b0),                                                                               // (terminated)
		.csr_write         (1'b0),                                                                               // (terminated)
		.csr_readdata      (),                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                               // (terminated)
		.almost_full_data  (),                                                                                   // (terminated)
		.almost_empty_data (),                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                               // (terminated)
		.out_empty         (),                                                                                   // (terminated)
		.in_error          (1'b0),                                                                               // (terminated)
		.out_error         (),                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                               // (terminated)
		.out_channel       ()                                                                                    // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (77),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (57),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (58),
		.PKT_TRANS_POSTED          (59),
		.PKT_TRANS_WRITE           (60),
		.PKT_TRANS_READ            (61),
		.PKT_TRANS_LOCK            (62),
		.PKT_SRC_ID_H              (85),
		.PKT_SRC_ID_L              (79),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (86),
		.PKT_BURSTWRAP_H           (69),
		.PKT_BURSTWRAP_L           (67),
		.PKT_BYTE_CNT_H            (66),
		.PKT_BYTE_CNT_L            (64),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (72),
		.PKT_BURST_SIZE_L          (70),
		.ST_CHANNEL_W              (99),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) ch4_yn1_l_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                           //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                //       clk_reset.reset
		.m0_address              (ch4_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ch4_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ch4_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ch4_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ch4_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ch4_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ch4_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ch4_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ch4_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ch4_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ch4_yn1_l_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ch4_yn1_l_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ch4_yn1_l_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ch4_yn1_l_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ch4_yn1_l_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ch4_yn1_l_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src90_ready),                                                    //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src90_valid),                                                    //                .valid
		.cp_data                 (cmd_xbar_demux_001_src90_data),                                                     //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src90_startofpacket),                                            //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src90_endofpacket),                                              //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src90_channel),                                                  //                .channel
		.rf_sink_ready           (ch4_yn1_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ch4_yn1_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ch4_yn1_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ch4_yn1_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ch4_yn1_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ch4_yn1_l_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ch4_yn1_l_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ch4_yn1_l_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ch4_yn1_l_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ch4_yn1_l_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ch4_yn1_l_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ch4_yn1_l_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (ch4_yn1_l_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (ch4_yn1_l_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ch4_yn1_l_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ch4_yn1_l_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                             //     (terminated)
		.m0_writeresponserequest (),                                                                                  //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                               //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ch4_yn1_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                           //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                // clk_reset.reset
		.in_data           (ch4_yn1_l_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ch4_yn1_l_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ch4_yn1_l_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ch4_yn1_l_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ch4_yn1_l_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ch4_yn1_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ch4_yn1_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ch4_yn1_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ch4_yn1_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ch4_yn1_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                             // (terminated)
		.csr_read          (1'b0),                                                                              // (terminated)
		.csr_write         (1'b0),                                                                              // (terminated)
		.csr_readdata      (),                                                                                  // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                              // (terminated)
		.almost_full_data  (),                                                                                  // (terminated)
		.almost_empty_data (),                                                                                  // (terminated)
		.in_empty          (1'b0),                                                                              // (terminated)
		.out_empty         (),                                                                                  // (terminated)
		.in_error          (1'b0),                                                                              // (terminated)
		.out_error         (),                                                                                  // (terminated)
		.in_channel        (1'b0),                                                                              // (terminated)
		.out_channel       ()                                                                                   // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (77),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (57),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (58),
		.PKT_TRANS_POSTED          (59),
		.PKT_TRANS_WRITE           (60),
		.PKT_TRANS_READ            (61),
		.PKT_TRANS_LOCK            (62),
		.PKT_SRC_ID_H              (85),
		.PKT_SRC_ID_L              (79),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (86),
		.PKT_BURSTWRAP_H           (69),
		.PKT_BURSTWRAP_L           (67),
		.PKT_BYTE_CNT_H            (66),
		.PKT_BYTE_CNT_L            (64),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (72),
		.PKT_BURST_SIZE_L          (70),
		.ST_CHANNEL_W              (99),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) ch4_yn2_u_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                           //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                //       clk_reset.reset
		.m0_address              (ch4_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ch4_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ch4_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ch4_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ch4_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ch4_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ch4_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ch4_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ch4_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ch4_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ch4_yn2_u_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ch4_yn2_u_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ch4_yn2_u_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ch4_yn2_u_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ch4_yn2_u_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ch4_yn2_u_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src91_ready),                                                    //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src91_valid),                                                    //                .valid
		.cp_data                 (cmd_xbar_demux_001_src91_data),                                                     //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src91_startofpacket),                                            //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src91_endofpacket),                                              //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src91_channel),                                                  //                .channel
		.rf_sink_ready           (ch4_yn2_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ch4_yn2_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ch4_yn2_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ch4_yn2_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ch4_yn2_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ch4_yn2_u_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ch4_yn2_u_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ch4_yn2_u_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ch4_yn2_u_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ch4_yn2_u_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ch4_yn2_u_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ch4_yn2_u_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (ch4_yn2_u_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (ch4_yn2_u_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ch4_yn2_u_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ch4_yn2_u_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                             //     (terminated)
		.m0_writeresponserequest (),                                                                                  //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                               //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ch4_yn2_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                           //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                // clk_reset.reset
		.in_data           (ch4_yn2_u_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ch4_yn2_u_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ch4_yn2_u_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ch4_yn2_u_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ch4_yn2_u_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ch4_yn2_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ch4_yn2_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ch4_yn2_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ch4_yn2_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ch4_yn2_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                             // (terminated)
		.csr_read          (1'b0),                                                                              // (terminated)
		.csr_write         (1'b0),                                                                              // (terminated)
		.csr_readdata      (),                                                                                  // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                              // (terminated)
		.almost_full_data  (),                                                                                  // (terminated)
		.almost_empty_data (),                                                                                  // (terminated)
		.in_empty          (1'b0),                                                                              // (terminated)
		.out_empty         (),                                                                                  // (terminated)
		.in_error          (1'b0),                                                                              // (terminated)
		.out_error         (),                                                                                  // (terminated)
		.in_channel        (1'b0),                                                                              // (terminated)
		.out_channel       ()                                                                                   // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (77),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (57),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (58),
		.PKT_TRANS_POSTED          (59),
		.PKT_TRANS_WRITE           (60),
		.PKT_TRANS_READ            (61),
		.PKT_TRANS_LOCK            (62),
		.PKT_SRC_ID_H              (85),
		.PKT_SRC_ID_L              (79),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (86),
		.PKT_BURSTWRAP_H           (69),
		.PKT_BURSTWRAP_L           (67),
		.PKT_BYTE_CNT_H            (66),
		.PKT_BYTE_CNT_L            (64),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (72),
		.PKT_BURST_SIZE_L          (70),
		.ST_CHANNEL_W              (99),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) ch4_yn2_mu_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                            //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                 //       clk_reset.reset
		.m0_address              (ch4_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ch4_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ch4_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ch4_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ch4_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ch4_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ch4_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ch4_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ch4_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ch4_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ch4_yn2_mu_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ch4_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ch4_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ch4_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ch4_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ch4_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src92_ready),                                                     //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src92_valid),                                                     //                .valid
		.cp_data                 (cmd_xbar_demux_001_src92_data),                                                      //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src92_startofpacket),                                             //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src92_endofpacket),                                               //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src92_channel),                                                   //                .channel
		.rf_sink_ready           (ch4_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ch4_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ch4_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ch4_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ch4_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ch4_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ch4_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ch4_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ch4_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ch4_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ch4_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ch4_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (ch4_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (ch4_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ch4_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ch4_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                              //     (terminated)
		.m0_writeresponserequest (),                                                                                   //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ch4_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                            //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                 // clk_reset.reset
		.in_data           (ch4_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ch4_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ch4_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ch4_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ch4_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ch4_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ch4_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ch4_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ch4_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ch4_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                              // (terminated)
		.csr_read          (1'b0),                                                                               // (terminated)
		.csr_write         (1'b0),                                                                               // (terminated)
		.csr_readdata      (),                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                               // (terminated)
		.almost_full_data  (),                                                                                   // (terminated)
		.almost_empty_data (),                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                               // (terminated)
		.out_empty         (),                                                                                   // (terminated)
		.in_error          (1'b0),                                                                               // (terminated)
		.out_error         (),                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                               // (terminated)
		.out_channel       ()                                                                                    // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (77),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (57),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (58),
		.PKT_TRANS_POSTED          (59),
		.PKT_TRANS_WRITE           (60),
		.PKT_TRANS_READ            (61),
		.PKT_TRANS_LOCK            (62),
		.PKT_SRC_ID_H              (85),
		.PKT_SRC_ID_L              (79),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (86),
		.PKT_BURSTWRAP_H           (69),
		.PKT_BURSTWRAP_L           (67),
		.PKT_BYTE_CNT_H            (66),
		.PKT_BYTE_CNT_L            (64),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (72),
		.PKT_BURST_SIZE_L          (70),
		.ST_CHANNEL_W              (99),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) ch4_yn2_ml_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                            //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                 //       clk_reset.reset
		.m0_address              (ch4_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ch4_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ch4_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ch4_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ch4_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ch4_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ch4_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ch4_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ch4_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ch4_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ch4_yn2_ml_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ch4_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ch4_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ch4_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ch4_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ch4_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src93_ready),                                                     //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src93_valid),                                                     //                .valid
		.cp_data                 (cmd_xbar_demux_001_src93_data),                                                      //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src93_startofpacket),                                             //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src93_endofpacket),                                               //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src93_channel),                                                   //                .channel
		.rf_sink_ready           (ch4_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ch4_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ch4_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ch4_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ch4_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ch4_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ch4_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ch4_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ch4_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ch4_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ch4_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ch4_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (ch4_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (ch4_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ch4_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ch4_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                              //     (terminated)
		.m0_writeresponserequest (),                                                                                   //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ch4_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                            //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                 // clk_reset.reset
		.in_data           (ch4_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ch4_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ch4_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ch4_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ch4_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ch4_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ch4_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ch4_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ch4_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ch4_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                              // (terminated)
		.csr_read          (1'b0),                                                                               // (terminated)
		.csr_write         (1'b0),                                                                               // (terminated)
		.csr_readdata      (),                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                               // (terminated)
		.almost_full_data  (),                                                                                   // (terminated)
		.almost_empty_data (),                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                               // (terminated)
		.out_empty         (),                                                                                   // (terminated)
		.in_error          (1'b0),                                                                               // (terminated)
		.out_error         (),                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                               // (terminated)
		.out_channel       ()                                                                                    // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (77),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (57),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (58),
		.PKT_TRANS_POSTED          (59),
		.PKT_TRANS_WRITE           (60),
		.PKT_TRANS_READ            (61),
		.PKT_TRANS_LOCK            (62),
		.PKT_SRC_ID_H              (85),
		.PKT_SRC_ID_L              (79),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (86),
		.PKT_BURSTWRAP_H           (69),
		.PKT_BURSTWRAP_L           (67),
		.PKT_BYTE_CNT_H            (66),
		.PKT_BYTE_CNT_L            (64),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (72),
		.PKT_BURST_SIZE_L          (70),
		.ST_CHANNEL_W              (99),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) ch4_yn2_l_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                           //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                //       clk_reset.reset
		.m0_address              (ch4_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ch4_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ch4_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ch4_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ch4_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ch4_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ch4_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ch4_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ch4_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ch4_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ch4_yn2_l_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ch4_yn2_l_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ch4_yn2_l_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ch4_yn2_l_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ch4_yn2_l_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ch4_yn2_l_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src94_ready),                                                    //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src94_valid),                                                    //                .valid
		.cp_data                 (cmd_xbar_demux_001_src94_data),                                                     //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src94_startofpacket),                                            //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src94_endofpacket),                                              //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src94_channel),                                                  //                .channel
		.rf_sink_ready           (ch4_yn2_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ch4_yn2_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ch4_yn2_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ch4_yn2_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ch4_yn2_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ch4_yn2_l_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ch4_yn2_l_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ch4_yn2_l_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ch4_yn2_l_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ch4_yn2_l_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ch4_yn2_l_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ch4_yn2_l_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (ch4_yn2_l_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (ch4_yn2_l_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ch4_yn2_l_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ch4_yn2_l_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                             //     (terminated)
		.m0_writeresponserequest (),                                                                                  //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                               //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ch4_yn2_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                           //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                // clk_reset.reset
		.in_data           (ch4_yn2_l_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ch4_yn2_l_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ch4_yn2_l_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ch4_yn2_l_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ch4_yn2_l_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ch4_yn2_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ch4_yn2_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ch4_yn2_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ch4_yn2_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ch4_yn2_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                             // (terminated)
		.csr_read          (1'b0),                                                                              // (terminated)
		.csr_write         (1'b0),                                                                              // (terminated)
		.csr_readdata      (),                                                                                  // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                              // (terminated)
		.almost_full_data  (),                                                                                  // (terminated)
		.almost_empty_data (),                                                                                  // (terminated)
		.in_empty          (1'b0),                                                                              // (terminated)
		.out_empty         (),                                                                                  // (terminated)
		.in_error          (1'b0),                                                                              // (terminated)
		.out_error         (),                                                                                  // (terminated)
		.in_channel        (1'b0),                                                                              // (terminated)
		.out_channel       ()                                                                                   // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (77),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (57),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (58),
		.PKT_TRANS_POSTED          (59),
		.PKT_TRANS_WRITE           (60),
		.PKT_TRANS_READ            (61),
		.PKT_TRANS_LOCK            (62),
		.PKT_SRC_ID_H              (85),
		.PKT_SRC_ID_L              (79),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (86),
		.PKT_BURSTWRAP_H           (69),
		.PKT_BURSTWRAP_L           (67),
		.PKT_BYTE_CNT_H            (66),
		.PKT_BYTE_CNT_L            (64),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (72),
		.PKT_BURST_SIZE_L          (70),
		.ST_CHANNEL_W              (99),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) ch4_yn3_u_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                           //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                //       clk_reset.reset
		.m0_address              (ch4_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ch4_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ch4_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ch4_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ch4_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ch4_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ch4_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ch4_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ch4_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ch4_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ch4_yn3_u_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ch4_yn3_u_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ch4_yn3_u_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ch4_yn3_u_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ch4_yn3_u_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ch4_yn3_u_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src95_ready),                                                    //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src95_valid),                                                    //                .valid
		.cp_data                 (cmd_xbar_demux_001_src95_data),                                                     //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src95_startofpacket),                                            //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src95_endofpacket),                                              //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src95_channel),                                                  //                .channel
		.rf_sink_ready           (ch4_yn3_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ch4_yn3_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ch4_yn3_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ch4_yn3_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ch4_yn3_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ch4_yn3_u_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ch4_yn3_u_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ch4_yn3_u_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ch4_yn3_u_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ch4_yn3_u_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ch4_yn3_u_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ch4_yn3_u_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (ch4_yn3_u_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (ch4_yn3_u_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ch4_yn3_u_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ch4_yn3_u_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                             //     (terminated)
		.m0_writeresponserequest (),                                                                                  //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                               //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ch4_yn3_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                           //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                // clk_reset.reset
		.in_data           (ch4_yn3_u_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ch4_yn3_u_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ch4_yn3_u_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ch4_yn3_u_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ch4_yn3_u_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ch4_yn3_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ch4_yn3_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ch4_yn3_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ch4_yn3_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ch4_yn3_u_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                             // (terminated)
		.csr_read          (1'b0),                                                                              // (terminated)
		.csr_write         (1'b0),                                                                              // (terminated)
		.csr_readdata      (),                                                                                  // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                              // (terminated)
		.almost_full_data  (),                                                                                  // (terminated)
		.almost_empty_data (),                                                                                  // (terminated)
		.in_empty          (1'b0),                                                                              // (terminated)
		.out_empty         (),                                                                                  // (terminated)
		.in_error          (1'b0),                                                                              // (terminated)
		.out_error         (),                                                                                  // (terminated)
		.in_channel        (1'b0),                                                                              // (terminated)
		.out_channel       ()                                                                                   // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (77),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (57),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (58),
		.PKT_TRANS_POSTED          (59),
		.PKT_TRANS_WRITE           (60),
		.PKT_TRANS_READ            (61),
		.PKT_TRANS_LOCK            (62),
		.PKT_SRC_ID_H              (85),
		.PKT_SRC_ID_L              (79),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (86),
		.PKT_BURSTWRAP_H           (69),
		.PKT_BURSTWRAP_L           (67),
		.PKT_BYTE_CNT_H            (66),
		.PKT_BYTE_CNT_L            (64),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (72),
		.PKT_BURST_SIZE_L          (70),
		.ST_CHANNEL_W              (99),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) ch4_yn3_mu_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                            //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                 //       clk_reset.reset
		.m0_address              (ch4_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ch4_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ch4_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ch4_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ch4_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ch4_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ch4_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ch4_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ch4_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ch4_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ch4_yn3_mu_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ch4_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ch4_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ch4_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ch4_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ch4_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src96_ready),                                                     //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src96_valid),                                                     //                .valid
		.cp_data                 (cmd_xbar_demux_001_src96_data),                                                      //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src96_startofpacket),                                             //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src96_endofpacket),                                               //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src96_channel),                                                   //                .channel
		.rf_sink_ready           (ch4_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ch4_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ch4_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ch4_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ch4_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ch4_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ch4_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ch4_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ch4_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ch4_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ch4_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ch4_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (ch4_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (ch4_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ch4_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ch4_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                              //     (terminated)
		.m0_writeresponserequest (),                                                                                   //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ch4_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                            //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                 // clk_reset.reset
		.in_data           (ch4_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ch4_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ch4_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ch4_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ch4_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ch4_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ch4_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ch4_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ch4_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ch4_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                              // (terminated)
		.csr_read          (1'b0),                                                                               // (terminated)
		.csr_write         (1'b0),                                                                               // (terminated)
		.csr_readdata      (),                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                               // (terminated)
		.almost_full_data  (),                                                                                   // (terminated)
		.almost_empty_data (),                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                               // (terminated)
		.out_empty         (),                                                                                   // (terminated)
		.in_error          (1'b0),                                                                               // (terminated)
		.out_error         (),                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                               // (terminated)
		.out_channel       ()                                                                                    // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (77),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (57),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (58),
		.PKT_TRANS_POSTED          (59),
		.PKT_TRANS_WRITE           (60),
		.PKT_TRANS_READ            (61),
		.PKT_TRANS_LOCK            (62),
		.PKT_SRC_ID_H              (85),
		.PKT_SRC_ID_L              (79),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (86),
		.PKT_BURSTWRAP_H           (69),
		.PKT_BURSTWRAP_L           (67),
		.PKT_BYTE_CNT_H            (66),
		.PKT_BYTE_CNT_L            (64),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (72),
		.PKT_BURST_SIZE_L          (70),
		.ST_CHANNEL_W              (99),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) ch4_yn3_ml_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                            //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                 //       clk_reset.reset
		.m0_address              (ch4_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ch4_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ch4_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ch4_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ch4_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ch4_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ch4_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ch4_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ch4_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ch4_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ch4_yn3_ml_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ch4_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ch4_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ch4_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ch4_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ch4_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src97_ready),                                                     //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src97_valid),                                                     //                .valid
		.cp_data                 (cmd_xbar_demux_001_src97_data),                                                      //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src97_startofpacket),                                             //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src97_endofpacket),                                               //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src97_channel),                                                   //                .channel
		.rf_sink_ready           (ch4_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ch4_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ch4_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ch4_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ch4_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ch4_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ch4_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ch4_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ch4_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ch4_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ch4_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ch4_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (ch4_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (ch4_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ch4_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ch4_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                              //     (terminated)
		.m0_writeresponserequest (),                                                                                   //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ch4_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                            //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                 // clk_reset.reset
		.in_data           (ch4_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ch4_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ch4_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ch4_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ch4_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ch4_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ch4_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ch4_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ch4_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ch4_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                              // (terminated)
		.csr_read          (1'b0),                                                                               // (terminated)
		.csr_write         (1'b0),                                                                               // (terminated)
		.csr_readdata      (),                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                               // (terminated)
		.almost_full_data  (),                                                                                   // (terminated)
		.almost_empty_data (),                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                               // (terminated)
		.out_empty         (),                                                                                   // (terminated)
		.in_error          (1'b0),                                                                               // (terminated)
		.out_error         (),                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                               // (terminated)
		.out_channel       ()                                                                                    // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (77),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (57),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (58),
		.PKT_TRANS_POSTED          (59),
		.PKT_TRANS_WRITE           (60),
		.PKT_TRANS_READ            (61),
		.PKT_TRANS_LOCK            (62),
		.PKT_SRC_ID_H              (85),
		.PKT_SRC_ID_L              (79),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (86),
		.PKT_BURSTWRAP_H           (69),
		.PKT_BURSTWRAP_L           (67),
		.PKT_BYTE_CNT_H            (66),
		.PKT_BYTE_CNT_L            (64),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (72),
		.PKT_BURST_SIZE_L          (70),
		.ST_CHANNEL_W              (99),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) ch4_yn3_l_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                           //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                //       clk_reset.reset
		.m0_address              (ch4_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ch4_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ch4_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ch4_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ch4_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ch4_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ch4_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ch4_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ch4_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ch4_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ch4_yn3_l_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ch4_yn3_l_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ch4_yn3_l_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ch4_yn3_l_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ch4_yn3_l_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ch4_yn3_l_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src98_ready),                                                    //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src98_valid),                                                    //                .valid
		.cp_data                 (cmd_xbar_demux_001_src98_data),                                                     //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src98_startofpacket),                                            //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src98_endofpacket),                                              //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src98_channel),                                                  //                .channel
		.rf_sink_ready           (ch4_yn3_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ch4_yn3_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ch4_yn3_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ch4_yn3_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ch4_yn3_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ch4_yn3_l_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ch4_yn3_l_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ch4_yn3_l_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ch4_yn3_l_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ch4_yn3_l_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ch4_yn3_l_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ch4_yn3_l_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (ch4_yn3_l_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (ch4_yn3_l_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ch4_yn3_l_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ch4_yn3_l_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                             //     (terminated)
		.m0_writeresponserequest (),                                                                                  //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                               //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ch4_yn3_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                           //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                // clk_reset.reset
		.in_data           (ch4_yn3_l_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ch4_yn3_l_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ch4_yn3_l_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ch4_yn3_l_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ch4_yn3_l_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ch4_yn3_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ch4_yn3_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ch4_yn3_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ch4_yn3_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ch4_yn3_l_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                             // (terminated)
		.csr_read          (1'b0),                                                                              // (terminated)
		.csr_write         (1'b0),                                                                              // (terminated)
		.csr_readdata      (),                                                                                  // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                              // (terminated)
		.almost_full_data  (),                                                                                  // (terminated)
		.almost_empty_data (),                                                                                  // (terminated)
		.in_empty          (1'b0),                                                                              // (terminated)
		.out_empty         (),                                                                                  // (terminated)
		.in_error          (1'b0),                                                                              // (terminated)
		.out_error         (),                                                                                  // (terminated)
		.in_channel        (1'b0),                                                                              // (terminated)
		.out_channel       ()                                                                                   // (terminated)
	);

	NIOS_SYSTEMV3_addr_router addr_router (
		.sink_ready         (nios_cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (nios_cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (nios_cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (nios_cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (nios_cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                                 //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                          // clk_reset.reset
		.src_ready          (addr_router_src_ready),                                                                   //       src.ready
		.src_valid          (addr_router_src_valid),                                                                   //          .valid
		.src_data           (addr_router_src_data),                                                                    //          .data
		.src_channel        (addr_router_src_channel),                                                                 //          .channel
		.src_startofpacket  (addr_router_src_startofpacket),                                                           //          .startofpacket
		.src_endofpacket    (addr_router_src_endofpacket)                                                              //          .endofpacket
	);

	NIOS_SYSTEMV3_addr_router_001 addr_router_001 (
		.sink_ready         (nios_cpu_data_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (nios_cpu_data_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (nios_cpu_data_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (nios_cpu_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (nios_cpu_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                          //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                   // clk_reset.reset
		.src_ready          (addr_router_001_src_ready),                                                        //       src.ready
		.src_valid          (addr_router_001_src_valid),                                                        //          .valid
		.src_data           (addr_router_001_src_data),                                                         //          .data
		.src_channel        (addr_router_001_src_channel),                                                      //          .channel
		.src_startofpacket  (addr_router_001_src_startofpacket),                                                //          .startofpacket
		.src_endofpacket    (addr_router_001_src_endofpacket)                                                   //          .endofpacket
	);

	NIOS_SYSTEMV3_id_router id_router (
		.sink_ready         (nios_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (nios_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (nios_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (nios_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (nios_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                        // clk_reset.reset
		.src_ready          (id_router_src_ready),                                                                   //       src.ready
		.src_valid          (id_router_src_valid),                                                                   //          .valid
		.src_data           (id_router_src_data),                                                                    //          .data
		.src_channel        (id_router_src_channel),                                                                 //          .channel
		.src_startofpacket  (id_router_src_startofpacket),                                                           //          .startofpacket
		.src_endofpacket    (id_router_src_endofpacket)                                                              //          .endofpacket
	);

	NIOS_SYSTEMV3_id_router id_router_001 (
		.sink_ready         (ram_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ram_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ram_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ram_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ram_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                           //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                // clk_reset.reset
		.src_ready          (id_router_001_src_ready),                                           //       src.ready
		.src_valid          (id_router_001_src_valid),                                           //          .valid
		.src_data           (id_router_001_src_data),                                            //          .data
		.src_channel        (id_router_001_src_channel),                                         //          .channel
		.src_startofpacket  (id_router_001_src_startofpacket),                                   //          .startofpacket
		.src_endofpacket    (id_router_001_src_endofpacket)                                      //          .endofpacket
	);

	NIOS_SYSTEMV3_id_router id_router_002 (
		.sink_ready         (ssram_uas_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ssram_uas_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ssram_uas_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ssram_uas_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ssram_uas_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                              //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                   // clk_reset.reset
		.src_ready          (id_router_002_src_ready),                                              //       src.ready
		.src_valid          (id_router_002_src_valid),                                              //          .valid
		.src_data           (id_router_002_src_data),                                               //          .data
		.src_channel        (id_router_002_src_channel),                                            //          .channel
		.src_startofpacket  (id_router_002_src_startofpacket),                                      //          .startofpacket
		.src_endofpacket    (id_router_002_src_endofpacket)                                         //          .endofpacket
	);

	NIOS_SYSTEMV3_id_router_003 id_router_003 (
		.sink_ready         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                                //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                                     // clk_reset.reset
		.src_ready          (id_router_003_src_ready),                                                                //       src.ready
		.src_valid          (id_router_003_src_valid),                                                                //          .valid
		.src_data           (id_router_003_src_data),                                                                 //          .data
		.src_channel        (id_router_003_src_channel),                                                              //          .channel
		.src_startofpacket  (id_router_003_src_startofpacket),                                                        //          .startofpacket
		.src_endofpacket    (id_router_003_src_endofpacket)                                                           //          .endofpacket
	);

	NIOS_SYSTEMV3_id_router_003 id_router_004 (
		.sink_ready         (lcd_control_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (lcd_control_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (lcd_control_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (lcd_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (lcd_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                      //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                           // clk_reset.reset
		.src_ready          (id_router_004_src_ready),                                                      //       src.ready
		.src_valid          (id_router_004_src_valid),                                                      //          .valid
		.src_data           (id_router_004_src_data),                                                       //          .data
		.src_channel        (id_router_004_src_channel),                                                    //          .channel
		.src_startofpacket  (id_router_004_src_startofpacket),                                              //          .startofpacket
		.src_endofpacket    (id_router_004_src_endofpacket)                                                 //          .endofpacket
	);

	NIOS_SYSTEMV3_id_router_003 id_router_005 (
		.sink_ready         (adc_on_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (adc_on_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (adc_on_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (adc_on_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (adc_on_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                              //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                   // clk_reset.reset
		.src_ready          (id_router_005_src_ready),                                              //       src.ready
		.src_valid          (id_router_005_src_valid),                                              //          .valid
		.src_data           (id_router_005_src_data),                                               //          .data
		.src_channel        (id_router_005_src_channel),                                            //          .channel
		.src_startofpacket  (id_router_005_src_startofpacket),                                      //          .startofpacket
		.src_endofpacket    (id_router_005_src_endofpacket)                                         //          .endofpacket
	);

	NIOS_SYSTEMV3_id_router_003 id_router_006 (
		.sink_ready         (fifo_adc_data_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (fifo_adc_data_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (fifo_adc_data_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (fifo_adc_data_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (fifo_adc_data_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                     //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                          // clk_reset.reset
		.src_ready          (id_router_006_src_ready),                                                     //       src.ready
		.src_valid          (id_router_006_src_valid),                                                     //          .valid
		.src_data           (id_router_006_src_data),                                                      //          .data
		.src_channel        (id_router_006_src_channel),                                                   //          .channel
		.src_startofpacket  (id_router_006_src_startofpacket),                                             //          .startofpacket
		.src_endofpacket    (id_router_006_src_endofpacket)                                                //          .endofpacket
	);

	NIOS_SYSTEMV3_id_router_003 id_router_007 (
		.sink_ready         (fifo_adc_data_valid_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (fifo_adc_data_valid_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (fifo_adc_data_valid_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (fifo_adc_data_valid_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (fifo_adc_data_valid_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                           //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                                // clk_reset.reset
		.src_ready          (id_router_007_src_ready),                                                           //       src.ready
		.src_valid          (id_router_007_src_valid),                                                           //          .valid
		.src_data           (id_router_007_src_data),                                                            //          .data
		.src_channel        (id_router_007_src_channel),                                                         //          .channel
		.src_startofpacket  (id_router_007_src_startofpacket),                                                   //          .startofpacket
		.src_endofpacket    (id_router_007_src_endofpacket)                                                      //          .endofpacket
	);

	NIOS_SYSTEMV3_id_router_003 id_router_008 (
		.sink_ready         (fifo_rst_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (fifo_rst_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (fifo_rst_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (fifo_rst_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (fifo_rst_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                     // clk_reset.reset
		.src_ready          (id_router_008_src_ready),                                                //       src.ready
		.src_valid          (id_router_008_src_valid),                                                //          .valid
		.src_data           (id_router_008_src_data),                                                 //          .data
		.src_channel        (id_router_008_src_channel),                                              //          .channel
		.src_startofpacket  (id_router_008_src_startofpacket),                                        //          .startofpacket
		.src_endofpacket    (id_router_008_src_endofpacket)                                           //          .endofpacket
	);

	NIOS_SYSTEMV3_id_router_003 id_router_009 (
		.sink_ready         (subtractor_on_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (subtractor_on_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (subtractor_on_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (subtractor_on_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (subtractor_on_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                     //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                          // clk_reset.reset
		.src_ready          (id_router_009_src_ready),                                                     //       src.ready
		.src_valid          (id_router_009_src_valid),                                                     //          .valid
		.src_data           (id_router_009_src_data),                                                      //          .data
		.src_channel        (id_router_009_src_channel),                                                   //          .channel
		.src_startofpacket  (id_router_009_src_startofpacket),                                             //          .startofpacket
		.src_endofpacket    (id_router_009_src_endofpacket)                                                //          .endofpacket
	);

	NIOS_SYSTEMV3_id_router_003 id_router_010 (
		.sink_ready         (ch0_timer_rst_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ch0_timer_rst_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ch0_timer_rst_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ch0_timer_rst_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ch0_timer_rst_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                     //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                          // clk_reset.reset
		.src_ready          (id_router_010_src_ready),                                                     //       src.ready
		.src_valid          (id_router_010_src_valid),                                                     //          .valid
		.src_data           (id_router_010_src_data),                                                      //          .data
		.src_channel        (id_router_010_src_channel),                                                   //          .channel
		.src_startofpacket  (id_router_010_src_startofpacket),                                             //          .startofpacket
		.src_endofpacket    (id_router_010_src_endofpacket)                                                //          .endofpacket
	);

	NIOS_SYSTEMV3_id_router_003 id_router_011 (
		.sink_ready         (detector_on_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (detector_on_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (detector_on_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (detector_on_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (detector_on_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                   //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                        // clk_reset.reset
		.src_ready          (id_router_011_src_ready),                                                   //       src.ready
		.src_valid          (id_router_011_src_valid),                                                   //          .valid
		.src_data           (id_router_011_src_data),                                                    //          .data
		.src_channel        (id_router_011_src_channel),                                                 //          .channel
		.src_startofpacket  (id_router_011_src_startofpacket),                                           //          .startofpacket
		.src_endofpacket    (id_router_011_src_endofpacket)                                              //          .endofpacket
	);

	NIOS_SYSTEMV3_id_router_003 id_router_012 (
		.sink_ready         (menu_down_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (menu_down_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (menu_down_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (menu_down_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (menu_down_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                 //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                      // clk_reset.reset
		.src_ready          (id_router_012_src_ready),                                                 //       src.ready
		.src_valid          (id_router_012_src_valid),                                                 //          .valid
		.src_data           (id_router_012_src_data),                                                  //          .data
		.src_channel        (id_router_012_src_channel),                                               //          .channel
		.src_startofpacket  (id_router_012_src_startofpacket),                                         //          .startofpacket
		.src_endofpacket    (id_router_012_src_endofpacket)                                            //          .endofpacket
	);

	NIOS_SYSTEMV3_id_router_003 id_router_013 (
		.sink_ready         (menu_up_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (menu_up_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (menu_up_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (menu_up_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (menu_up_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                    // clk_reset.reset
		.src_ready          (id_router_013_src_ready),                                               //       src.ready
		.src_valid          (id_router_013_src_valid),                                               //          .valid
		.src_data           (id_router_013_src_data),                                                //          .data
		.src_channel        (id_router_013_src_channel),                                             //          .channel
		.src_startofpacket  (id_router_013_src_startofpacket),                                       //          .startofpacket
		.src_endofpacket    (id_router_013_src_endofpacket)                                          //          .endofpacket
	);

	NIOS_SYSTEMV3_id_router_003 id_router_014 (
		.sink_ready         (menu_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (menu_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (menu_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (menu_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (menu_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                            //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                 // clk_reset.reset
		.src_ready          (id_router_014_src_ready),                                            //       src.ready
		.src_valid          (id_router_014_src_valid),                                            //          .valid
		.src_data           (id_router_014_src_data),                                             //          .data
		.src_channel        (id_router_014_src_channel),                                          //          .channel
		.src_startofpacket  (id_router_014_src_startofpacket),                                    //          .startofpacket
		.src_endofpacket    (id_router_014_src_endofpacket)                                       //          .endofpacket
	);

	NIOS_SYSTEMV3_id_router_003 id_router_015 (
		.sink_ready         (ch0_thresh_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ch0_thresh_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ch0_thresh_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ch0_thresh_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ch0_thresh_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                  //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                       // clk_reset.reset
		.src_ready          (id_router_015_src_ready),                                                  //       src.ready
		.src_valid          (id_router_015_src_valid),                                                  //          .valid
		.src_data           (id_router_015_src_data),                                                   //          .data
		.src_channel        (id_router_015_src_channel),                                                //          .channel
		.src_startofpacket  (id_router_015_src_startofpacket),                                          //          .startofpacket
		.src_endofpacket    (id_router_015_src_endofpacket)                                             //          .endofpacket
	);

	NIOS_SYSTEMV3_id_router_003 id_router_016 (
		.sink_ready         (ch0_rd_peak_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ch0_rd_peak_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ch0_rd_peak_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ch0_rd_peak_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ch0_rd_peak_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                   //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                        // clk_reset.reset
		.src_ready          (id_router_016_src_ready),                                                   //       src.ready
		.src_valid          (id_router_016_src_valid),                                                   //          .valid
		.src_data           (id_router_016_src_data),                                                    //          .data
		.src_channel        (id_router_016_src_channel),                                                 //          .channel
		.src_startofpacket  (id_router_016_src_startofpacket),                                           //          .startofpacket
		.src_endofpacket    (id_router_016_src_endofpacket)                                              //          .endofpacket
	);

	NIOS_SYSTEMV3_id_router_003 id_router_017 (
		.sink_ready         (ch0_peak_found_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ch0_peak_found_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ch0_peak_found_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ch0_peak_found_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ch0_peak_found_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                      //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                           // clk_reset.reset
		.src_ready          (id_router_017_src_ready),                                                      //       src.ready
		.src_valid          (id_router_017_src_valid),                                                      //          .valid
		.src_data           (id_router_017_src_data),                                                       //          .data
		.src_channel        (id_router_017_src_channel),                                                    //          .channel
		.src_startofpacket  (id_router_017_src_startofpacket),                                              //          .startofpacket
		.src_endofpacket    (id_router_017_src_endofpacket)                                                 //          .endofpacket
	);

	NIOS_SYSTEMV3_id_router_003 id_router_018 (
		.sink_ready         (ch0_yn1_l_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ch0_yn1_l_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ch0_yn1_l_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ch0_yn1_l_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ch0_yn1_l_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                 //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                      // clk_reset.reset
		.src_ready          (id_router_018_src_ready),                                                 //       src.ready
		.src_valid          (id_router_018_src_valid),                                                 //          .valid
		.src_data           (id_router_018_src_data),                                                  //          .data
		.src_channel        (id_router_018_src_channel),                                               //          .channel
		.src_startofpacket  (id_router_018_src_startofpacket),                                         //          .startofpacket
		.src_endofpacket    (id_router_018_src_endofpacket)                                            //          .endofpacket
	);

	NIOS_SYSTEMV3_id_router_003 id_router_019 (
		.sink_ready         (ch0_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ch0_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ch0_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ch0_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ch0_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                  //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                       // clk_reset.reset
		.src_ready          (id_router_019_src_ready),                                                  //       src.ready
		.src_valid          (id_router_019_src_valid),                                                  //          .valid
		.src_data           (id_router_019_src_data),                                                   //          .data
		.src_channel        (id_router_019_src_channel),                                                //          .channel
		.src_startofpacket  (id_router_019_src_startofpacket),                                          //          .startofpacket
		.src_endofpacket    (id_router_019_src_endofpacket)                                             //          .endofpacket
	);

	NIOS_SYSTEMV3_id_router_003 id_router_020 (
		.sink_ready         (ch0_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ch0_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ch0_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ch0_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ch0_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                  //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                       // clk_reset.reset
		.src_ready          (id_router_020_src_ready),                                                  //       src.ready
		.src_valid          (id_router_020_src_valid),                                                  //          .valid
		.src_data           (id_router_020_src_data),                                                   //          .data
		.src_channel        (id_router_020_src_channel),                                                //          .channel
		.src_startofpacket  (id_router_020_src_startofpacket),                                          //          .startofpacket
		.src_endofpacket    (id_router_020_src_endofpacket)                                             //          .endofpacket
	);

	NIOS_SYSTEMV3_id_router_003 id_router_021 (
		.sink_ready         (ch0_yn1_u_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ch0_yn1_u_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ch0_yn1_u_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ch0_yn1_u_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ch0_yn1_u_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                 //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                      // clk_reset.reset
		.src_ready          (id_router_021_src_ready),                                                 //       src.ready
		.src_valid          (id_router_021_src_valid),                                                 //          .valid
		.src_data           (id_router_021_src_data),                                                  //          .data
		.src_channel        (id_router_021_src_channel),                                               //          .channel
		.src_startofpacket  (id_router_021_src_startofpacket),                                         //          .startofpacket
		.src_endofpacket    (id_router_021_src_endofpacket)                                            //          .endofpacket
	);

	NIOS_SYSTEMV3_id_router_003 id_router_022 (
		.sink_ready         (ch0_time_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ch0_time_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ch0_time_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ch0_time_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ch0_time_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                     // clk_reset.reset
		.src_ready          (id_router_022_src_ready),                                                //       src.ready
		.src_valid          (id_router_022_src_valid),                                                //          .valid
		.src_data           (id_router_022_src_data),                                                 //          .data
		.src_channel        (id_router_022_src_channel),                                              //          .channel
		.src_startofpacket  (id_router_022_src_startofpacket),                                        //          .startofpacket
		.src_endofpacket    (id_router_022_src_endofpacket)                                           //          .endofpacket
	);

	NIOS_SYSTEMV3_id_router_003 id_router_023 (
		.sink_ready         (ch0_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ch0_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ch0_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ch0_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ch0_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                  //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                       // clk_reset.reset
		.src_ready          (id_router_023_src_ready),                                                  //       src.ready
		.src_valid          (id_router_023_src_valid),                                                  //          .valid
		.src_data           (id_router_023_src_data),                                                   //          .data
		.src_channel        (id_router_023_src_channel),                                                //          .channel
		.src_startofpacket  (id_router_023_src_startofpacket),                                          //          .startofpacket
		.src_endofpacket    (id_router_023_src_endofpacket)                                             //          .endofpacket
	);

	NIOS_SYSTEMV3_id_router_003 id_router_024 (
		.sink_ready         (ch0_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ch0_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ch0_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ch0_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ch0_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                  //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                       // clk_reset.reset
		.src_ready          (id_router_024_src_ready),                                                  //       src.ready
		.src_valid          (id_router_024_src_valid),                                                  //          .valid
		.src_data           (id_router_024_src_data),                                                   //          .data
		.src_channel        (id_router_024_src_channel),                                                //          .channel
		.src_startofpacket  (id_router_024_src_startofpacket),                                          //          .startofpacket
		.src_endofpacket    (id_router_024_src_endofpacket)                                             //          .endofpacket
	);

	NIOS_SYSTEMV3_id_router_003 id_router_025 (
		.sink_ready         (ch0_yn2_u_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ch0_yn2_u_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ch0_yn2_u_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ch0_yn2_u_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ch0_yn2_u_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                 //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                      // clk_reset.reset
		.src_ready          (id_router_025_src_ready),                                                 //       src.ready
		.src_valid          (id_router_025_src_valid),                                                 //          .valid
		.src_data           (id_router_025_src_data),                                                  //          .data
		.src_channel        (id_router_025_src_channel),                                               //          .channel
		.src_startofpacket  (id_router_025_src_startofpacket),                                         //          .startofpacket
		.src_endofpacket    (id_router_025_src_endofpacket)                                            //          .endofpacket
	);

	NIOS_SYSTEMV3_id_router_003 id_router_026 (
		.sink_ready         (ch0_yn2_l_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ch0_yn2_l_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ch0_yn2_l_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ch0_yn2_l_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ch0_yn2_l_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                 //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                      // clk_reset.reset
		.src_ready          (id_router_026_src_ready),                                                 //       src.ready
		.src_valid          (id_router_026_src_valid),                                                 //          .valid
		.src_data           (id_router_026_src_data),                                                  //          .data
		.src_channel        (id_router_026_src_channel),                                               //          .channel
		.src_startofpacket  (id_router_026_src_startofpacket),                                         //          .startofpacket
		.src_endofpacket    (id_router_026_src_endofpacket)                                            //          .endofpacket
	);

	NIOS_SYSTEMV3_id_router_003 id_router_027 (
		.sink_ready         (ch0_yn3_l_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ch0_yn3_l_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ch0_yn3_l_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ch0_yn3_l_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ch0_yn3_l_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                 //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                      // clk_reset.reset
		.src_ready          (id_router_027_src_ready),                                                 //       src.ready
		.src_valid          (id_router_027_src_valid),                                                 //          .valid
		.src_data           (id_router_027_src_data),                                                  //          .data
		.src_channel        (id_router_027_src_channel),                                               //          .channel
		.src_startofpacket  (id_router_027_src_startofpacket),                                         //          .startofpacket
		.src_endofpacket    (id_router_027_src_endofpacket)                                            //          .endofpacket
	);

	NIOS_SYSTEMV3_id_router_003 id_router_028 (
		.sink_ready         (ch0_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ch0_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ch0_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ch0_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ch0_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                  //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                       // clk_reset.reset
		.src_ready          (id_router_028_src_ready),                                                  //       src.ready
		.src_valid          (id_router_028_src_valid),                                                  //          .valid
		.src_data           (id_router_028_src_data),                                                   //          .data
		.src_channel        (id_router_028_src_channel),                                                //          .channel
		.src_startofpacket  (id_router_028_src_startofpacket),                                          //          .startofpacket
		.src_endofpacket    (id_router_028_src_endofpacket)                                             //          .endofpacket
	);

	NIOS_SYSTEMV3_id_router_003 id_router_029 (
		.sink_ready         (ch0_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ch0_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ch0_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ch0_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ch0_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                  //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                       // clk_reset.reset
		.src_ready          (id_router_029_src_ready),                                                  //       src.ready
		.src_valid          (id_router_029_src_valid),                                                  //          .valid
		.src_data           (id_router_029_src_data),                                                   //          .data
		.src_channel        (id_router_029_src_channel),                                                //          .channel
		.src_startofpacket  (id_router_029_src_startofpacket),                                          //          .startofpacket
		.src_endofpacket    (id_router_029_src_endofpacket)                                             //          .endofpacket
	);

	NIOS_SYSTEMV3_id_router_003 id_router_030 (
		.sink_ready         (ch0_yn3_u_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ch0_yn3_u_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ch0_yn3_u_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ch0_yn3_u_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ch0_yn3_u_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                 //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                      // clk_reset.reset
		.src_ready          (id_router_030_src_ready),                                                 //       src.ready
		.src_valid          (id_router_030_src_valid),                                                 //          .valid
		.src_data           (id_router_030_src_data),                                                  //          .data
		.src_channel        (id_router_030_src_channel),                                               //          .channel
		.src_startofpacket  (id_router_030_src_startofpacket),                                         //          .startofpacket
		.src_endofpacket    (id_router_030_src_endofpacket)                                            //          .endofpacket
	);

	NIOS_SYSTEMV3_id_router_003 id_router_031 (
		.sink_ready         (ch1_timer_rst_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ch1_timer_rst_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ch1_timer_rst_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ch1_timer_rst_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ch1_timer_rst_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                     //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                          // clk_reset.reset
		.src_ready          (id_router_031_src_ready),                                                     //       src.ready
		.src_valid          (id_router_031_src_valid),                                                     //          .valid
		.src_data           (id_router_031_src_data),                                                      //          .data
		.src_channel        (id_router_031_src_channel),                                                   //          .channel
		.src_startofpacket  (id_router_031_src_startofpacket),                                             //          .startofpacket
		.src_endofpacket    (id_router_031_src_endofpacket)                                                //          .endofpacket
	);

	NIOS_SYSTEMV3_id_router_003 id_router_032 (
		.sink_ready         (ch1_thresh_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ch1_thresh_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ch1_thresh_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ch1_thresh_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ch1_thresh_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                  //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                       // clk_reset.reset
		.src_ready          (id_router_032_src_ready),                                                  //       src.ready
		.src_valid          (id_router_032_src_valid),                                                  //          .valid
		.src_data           (id_router_032_src_data),                                                   //          .data
		.src_channel        (id_router_032_src_channel),                                                //          .channel
		.src_startofpacket  (id_router_032_src_startofpacket),                                          //          .startofpacket
		.src_endofpacket    (id_router_032_src_endofpacket)                                             //          .endofpacket
	);

	NIOS_SYSTEMV3_id_router_003 id_router_033 (
		.sink_ready         (ch1_rd_peak_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ch1_rd_peak_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ch1_rd_peak_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ch1_rd_peak_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ch1_rd_peak_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                   //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                        // clk_reset.reset
		.src_ready          (id_router_033_src_ready),                                                   //       src.ready
		.src_valid          (id_router_033_src_valid),                                                   //          .valid
		.src_data           (id_router_033_src_data),                                                    //          .data
		.src_channel        (id_router_033_src_channel),                                                 //          .channel
		.src_startofpacket  (id_router_033_src_startofpacket),                                           //          .startofpacket
		.src_endofpacket    (id_router_033_src_endofpacket)                                              //          .endofpacket
	);

	NIOS_SYSTEMV3_id_router_003 id_router_034 (
		.sink_ready         (ch1_peak_found_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ch1_peak_found_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ch1_peak_found_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ch1_peak_found_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ch1_peak_found_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                      //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                           // clk_reset.reset
		.src_ready          (id_router_034_src_ready),                                                      //       src.ready
		.src_valid          (id_router_034_src_valid),                                                      //          .valid
		.src_data           (id_router_034_src_data),                                                       //          .data
		.src_channel        (id_router_034_src_channel),                                                    //          .channel
		.src_startofpacket  (id_router_034_src_startofpacket),                                              //          .startofpacket
		.src_endofpacket    (id_router_034_src_endofpacket)                                                 //          .endofpacket
	);

	NIOS_SYSTEMV3_id_router_003 id_router_035 (
		.sink_ready         (ch1_time_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ch1_time_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ch1_time_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ch1_time_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ch1_time_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                     // clk_reset.reset
		.src_ready          (id_router_035_src_ready),                                                //       src.ready
		.src_valid          (id_router_035_src_valid),                                                //          .valid
		.src_data           (id_router_035_src_data),                                                 //          .data
		.src_channel        (id_router_035_src_channel),                                              //          .channel
		.src_startofpacket  (id_router_035_src_startofpacket),                                        //          .startofpacket
		.src_endofpacket    (id_router_035_src_endofpacket)                                           //          .endofpacket
	);

	NIOS_SYSTEMV3_id_router_003 id_router_036 (
		.sink_ready         (ch1_yn1_u_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ch1_yn1_u_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ch1_yn1_u_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ch1_yn1_u_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ch1_yn1_u_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                 //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                      // clk_reset.reset
		.src_ready          (id_router_036_src_ready),                                                 //       src.ready
		.src_valid          (id_router_036_src_valid),                                                 //          .valid
		.src_data           (id_router_036_src_data),                                                  //          .data
		.src_channel        (id_router_036_src_channel),                                               //          .channel
		.src_startofpacket  (id_router_036_src_startofpacket),                                         //          .startofpacket
		.src_endofpacket    (id_router_036_src_endofpacket)                                            //          .endofpacket
	);

	NIOS_SYSTEMV3_id_router_003 id_router_037 (
		.sink_ready         (ch1_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ch1_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ch1_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ch1_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ch1_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                  //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                       // clk_reset.reset
		.src_ready          (id_router_037_src_ready),                                                  //       src.ready
		.src_valid          (id_router_037_src_valid),                                                  //          .valid
		.src_data           (id_router_037_src_data),                                                   //          .data
		.src_channel        (id_router_037_src_channel),                                                //          .channel
		.src_startofpacket  (id_router_037_src_startofpacket),                                          //          .startofpacket
		.src_endofpacket    (id_router_037_src_endofpacket)                                             //          .endofpacket
	);

	NIOS_SYSTEMV3_id_router_003 id_router_038 (
		.sink_ready         (ch1_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ch1_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ch1_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ch1_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ch1_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                  //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                       // clk_reset.reset
		.src_ready          (id_router_038_src_ready),                                                  //       src.ready
		.src_valid          (id_router_038_src_valid),                                                  //          .valid
		.src_data           (id_router_038_src_data),                                                   //          .data
		.src_channel        (id_router_038_src_channel),                                                //          .channel
		.src_startofpacket  (id_router_038_src_startofpacket),                                          //          .startofpacket
		.src_endofpacket    (id_router_038_src_endofpacket)                                             //          .endofpacket
	);

	NIOS_SYSTEMV3_id_router_003 id_router_039 (
		.sink_ready         (ch1_yn1_l_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ch1_yn1_l_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ch1_yn1_l_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ch1_yn1_l_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ch1_yn1_l_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                 //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                      // clk_reset.reset
		.src_ready          (id_router_039_src_ready),                                                 //       src.ready
		.src_valid          (id_router_039_src_valid),                                                 //          .valid
		.src_data           (id_router_039_src_data),                                                  //          .data
		.src_channel        (id_router_039_src_channel),                                               //          .channel
		.src_startofpacket  (id_router_039_src_startofpacket),                                         //          .startofpacket
		.src_endofpacket    (id_router_039_src_endofpacket)                                            //          .endofpacket
	);

	NIOS_SYSTEMV3_id_router_003 id_router_040 (
		.sink_ready         (ch1_yn2_u_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ch1_yn2_u_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ch1_yn2_u_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ch1_yn2_u_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ch1_yn2_u_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                 //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                      // clk_reset.reset
		.src_ready          (id_router_040_src_ready),                                                 //       src.ready
		.src_valid          (id_router_040_src_valid),                                                 //          .valid
		.src_data           (id_router_040_src_data),                                                  //          .data
		.src_channel        (id_router_040_src_channel),                                               //          .channel
		.src_startofpacket  (id_router_040_src_startofpacket),                                         //          .startofpacket
		.src_endofpacket    (id_router_040_src_endofpacket)                                            //          .endofpacket
	);

	NIOS_SYSTEMV3_id_router_003 id_router_041 (
		.sink_ready         (ch1_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ch1_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ch1_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ch1_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ch1_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                  //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                       // clk_reset.reset
		.src_ready          (id_router_041_src_ready),                                                  //       src.ready
		.src_valid          (id_router_041_src_valid),                                                  //          .valid
		.src_data           (id_router_041_src_data),                                                   //          .data
		.src_channel        (id_router_041_src_channel),                                                //          .channel
		.src_startofpacket  (id_router_041_src_startofpacket),                                          //          .startofpacket
		.src_endofpacket    (id_router_041_src_endofpacket)                                             //          .endofpacket
	);

	NIOS_SYSTEMV3_id_router_003 id_router_042 (
		.sink_ready         (ch1_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ch1_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ch1_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ch1_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ch1_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                  //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                       // clk_reset.reset
		.src_ready          (id_router_042_src_ready),                                                  //       src.ready
		.src_valid          (id_router_042_src_valid),                                                  //          .valid
		.src_data           (id_router_042_src_data),                                                   //          .data
		.src_channel        (id_router_042_src_channel),                                                //          .channel
		.src_startofpacket  (id_router_042_src_startofpacket),                                          //          .startofpacket
		.src_endofpacket    (id_router_042_src_endofpacket)                                             //          .endofpacket
	);

	NIOS_SYSTEMV3_id_router_003 id_router_043 (
		.sink_ready         (ch1_yn2_l_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ch1_yn2_l_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ch1_yn2_l_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ch1_yn2_l_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ch1_yn2_l_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                 //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                      // clk_reset.reset
		.src_ready          (id_router_043_src_ready),                                                 //       src.ready
		.src_valid          (id_router_043_src_valid),                                                 //          .valid
		.src_data           (id_router_043_src_data),                                                  //          .data
		.src_channel        (id_router_043_src_channel),                                               //          .channel
		.src_startofpacket  (id_router_043_src_startofpacket),                                         //          .startofpacket
		.src_endofpacket    (id_router_043_src_endofpacket)                                            //          .endofpacket
	);

	NIOS_SYSTEMV3_id_router_003 id_router_044 (
		.sink_ready         (ch1_yn3_u_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ch1_yn3_u_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ch1_yn3_u_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ch1_yn3_u_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ch1_yn3_u_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                 //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                      // clk_reset.reset
		.src_ready          (id_router_044_src_ready),                                                 //       src.ready
		.src_valid          (id_router_044_src_valid),                                                 //          .valid
		.src_data           (id_router_044_src_data),                                                  //          .data
		.src_channel        (id_router_044_src_channel),                                               //          .channel
		.src_startofpacket  (id_router_044_src_startofpacket),                                         //          .startofpacket
		.src_endofpacket    (id_router_044_src_endofpacket)                                            //          .endofpacket
	);

	NIOS_SYSTEMV3_id_router_003 id_router_045 (
		.sink_ready         (ch1_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ch1_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ch1_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ch1_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ch1_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                  //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                       // clk_reset.reset
		.src_ready          (id_router_045_src_ready),                                                  //       src.ready
		.src_valid          (id_router_045_src_valid),                                                  //          .valid
		.src_data           (id_router_045_src_data),                                                   //          .data
		.src_channel        (id_router_045_src_channel),                                                //          .channel
		.src_startofpacket  (id_router_045_src_startofpacket),                                          //          .startofpacket
		.src_endofpacket    (id_router_045_src_endofpacket)                                             //          .endofpacket
	);

	NIOS_SYSTEMV3_id_router_003 id_router_046 (
		.sink_ready         (ch1_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ch1_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ch1_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ch1_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ch1_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                  //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                       // clk_reset.reset
		.src_ready          (id_router_046_src_ready),                                                  //       src.ready
		.src_valid          (id_router_046_src_valid),                                                  //          .valid
		.src_data           (id_router_046_src_data),                                                   //          .data
		.src_channel        (id_router_046_src_channel),                                                //          .channel
		.src_startofpacket  (id_router_046_src_startofpacket),                                          //          .startofpacket
		.src_endofpacket    (id_router_046_src_endofpacket)                                             //          .endofpacket
	);

	NIOS_SYSTEMV3_id_router_003 id_router_047 (
		.sink_ready         (ch1_yn3_l_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ch1_yn3_l_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ch1_yn3_l_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ch1_yn3_l_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ch1_yn3_l_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                 //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                      // clk_reset.reset
		.src_ready          (id_router_047_src_ready),                                                 //       src.ready
		.src_valid          (id_router_047_src_valid),                                                 //          .valid
		.src_data           (id_router_047_src_data),                                                  //          .data
		.src_channel        (id_router_047_src_channel),                                               //          .channel
		.src_startofpacket  (id_router_047_src_startofpacket),                                         //          .startofpacket
		.src_endofpacket    (id_router_047_src_endofpacket)                                            //          .endofpacket
	);

	NIOS_SYSTEMV3_id_router_003 id_router_048 (
		.sink_ready         (ch2_timer_rst_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ch2_timer_rst_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ch2_timer_rst_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ch2_timer_rst_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ch2_timer_rst_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                     //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                          // clk_reset.reset
		.src_ready          (id_router_048_src_ready),                                                     //       src.ready
		.src_valid          (id_router_048_src_valid),                                                     //          .valid
		.src_data           (id_router_048_src_data),                                                      //          .data
		.src_channel        (id_router_048_src_channel),                                                   //          .channel
		.src_startofpacket  (id_router_048_src_startofpacket),                                             //          .startofpacket
		.src_endofpacket    (id_router_048_src_endofpacket)                                                //          .endofpacket
	);

	NIOS_SYSTEMV3_id_router_003 id_router_049 (
		.sink_ready         (ch2_thresh_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ch2_thresh_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ch2_thresh_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ch2_thresh_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ch2_thresh_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                  //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                       // clk_reset.reset
		.src_ready          (id_router_049_src_ready),                                                  //       src.ready
		.src_valid          (id_router_049_src_valid),                                                  //          .valid
		.src_data           (id_router_049_src_data),                                                   //          .data
		.src_channel        (id_router_049_src_channel),                                                //          .channel
		.src_startofpacket  (id_router_049_src_startofpacket),                                          //          .startofpacket
		.src_endofpacket    (id_router_049_src_endofpacket)                                             //          .endofpacket
	);

	NIOS_SYSTEMV3_id_router_003 id_router_050 (
		.sink_ready         (ch2_rd_peak_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ch2_rd_peak_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ch2_rd_peak_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ch2_rd_peak_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ch2_rd_peak_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                   //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                        // clk_reset.reset
		.src_ready          (id_router_050_src_ready),                                                   //       src.ready
		.src_valid          (id_router_050_src_valid),                                                   //          .valid
		.src_data           (id_router_050_src_data),                                                    //          .data
		.src_channel        (id_router_050_src_channel),                                                 //          .channel
		.src_startofpacket  (id_router_050_src_startofpacket),                                           //          .startofpacket
		.src_endofpacket    (id_router_050_src_endofpacket)                                              //          .endofpacket
	);

	NIOS_SYSTEMV3_id_router_003 id_router_051 (
		.sink_ready         (ch2_peak_found_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ch2_peak_found_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ch2_peak_found_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ch2_peak_found_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ch2_peak_found_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                      //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                           // clk_reset.reset
		.src_ready          (id_router_051_src_ready),                                                      //       src.ready
		.src_valid          (id_router_051_src_valid),                                                      //          .valid
		.src_data           (id_router_051_src_data),                                                       //          .data
		.src_channel        (id_router_051_src_channel),                                                    //          .channel
		.src_startofpacket  (id_router_051_src_startofpacket),                                              //          .startofpacket
		.src_endofpacket    (id_router_051_src_endofpacket)                                                 //          .endofpacket
	);

	NIOS_SYSTEMV3_id_router_003 id_router_052 (
		.sink_ready         (ch2_time_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ch2_time_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ch2_time_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ch2_time_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ch2_time_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                     // clk_reset.reset
		.src_ready          (id_router_052_src_ready),                                                //       src.ready
		.src_valid          (id_router_052_src_valid),                                                //          .valid
		.src_data           (id_router_052_src_data),                                                 //          .data
		.src_channel        (id_router_052_src_channel),                                              //          .channel
		.src_startofpacket  (id_router_052_src_startofpacket),                                        //          .startofpacket
		.src_endofpacket    (id_router_052_src_endofpacket)                                           //          .endofpacket
	);

	NIOS_SYSTEMV3_id_router_003 id_router_053 (
		.sink_ready         (ch2_yn1_u_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ch2_yn1_u_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ch2_yn1_u_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ch2_yn1_u_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ch2_yn1_u_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                 //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                      // clk_reset.reset
		.src_ready          (id_router_053_src_ready),                                                 //       src.ready
		.src_valid          (id_router_053_src_valid),                                                 //          .valid
		.src_data           (id_router_053_src_data),                                                  //          .data
		.src_channel        (id_router_053_src_channel),                                               //          .channel
		.src_startofpacket  (id_router_053_src_startofpacket),                                         //          .startofpacket
		.src_endofpacket    (id_router_053_src_endofpacket)                                            //          .endofpacket
	);

	NIOS_SYSTEMV3_id_router_003 id_router_054 (
		.sink_ready         (ch2_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ch2_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ch2_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ch2_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ch2_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                  //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                       // clk_reset.reset
		.src_ready          (id_router_054_src_ready),                                                  //       src.ready
		.src_valid          (id_router_054_src_valid),                                                  //          .valid
		.src_data           (id_router_054_src_data),                                                   //          .data
		.src_channel        (id_router_054_src_channel),                                                //          .channel
		.src_startofpacket  (id_router_054_src_startofpacket),                                          //          .startofpacket
		.src_endofpacket    (id_router_054_src_endofpacket)                                             //          .endofpacket
	);

	NIOS_SYSTEMV3_id_router_003 id_router_055 (
		.sink_ready         (ch2_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ch2_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ch2_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ch2_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ch2_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                  //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                       // clk_reset.reset
		.src_ready          (id_router_055_src_ready),                                                  //       src.ready
		.src_valid          (id_router_055_src_valid),                                                  //          .valid
		.src_data           (id_router_055_src_data),                                                   //          .data
		.src_channel        (id_router_055_src_channel),                                                //          .channel
		.src_startofpacket  (id_router_055_src_startofpacket),                                          //          .startofpacket
		.src_endofpacket    (id_router_055_src_endofpacket)                                             //          .endofpacket
	);

	NIOS_SYSTEMV3_id_router_003 id_router_056 (
		.sink_ready         (ch2_yn1_l_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ch2_yn1_l_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ch2_yn1_l_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ch2_yn1_l_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ch2_yn1_l_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                 //       clk.clk
		.reset              (nios_cpu_jtag_debug_module_reset_reset),                                  // clk_reset.reset
		.src_ready          (id_router_056_src_ready),                                                 //       src.ready
		.src_valid          (id_router_056_src_valid),                                                 //          .valid
		.src_data           (id_router_056_src_data),                                                  //          .data
		.src_channel        (id_router_056_src_channel),                                               //          .channel
		.src_startofpacket  (id_router_056_src_startofpacket),                                         //          .startofpacket
		.src_endofpacket    (id_router_056_src_endofpacket)                                            //          .endofpacket
	);

	NIOS_SYSTEMV3_id_router_003 id_router_057 (
		.sink_ready         (ch2_yn2_u_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ch2_yn2_u_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ch2_yn2_u_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ch2_yn2_u_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ch2_yn2_u_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                 //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                      // clk_reset.reset
		.src_ready          (id_router_057_src_ready),                                                 //       src.ready
		.src_valid          (id_router_057_src_valid),                                                 //          .valid
		.src_data           (id_router_057_src_data),                                                  //          .data
		.src_channel        (id_router_057_src_channel),                                               //          .channel
		.src_startofpacket  (id_router_057_src_startofpacket),                                         //          .startofpacket
		.src_endofpacket    (id_router_057_src_endofpacket)                                            //          .endofpacket
	);

	NIOS_SYSTEMV3_id_router_003 id_router_058 (
		.sink_ready         (ch2_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ch2_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ch2_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ch2_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ch2_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                  //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                       // clk_reset.reset
		.src_ready          (id_router_058_src_ready),                                                  //       src.ready
		.src_valid          (id_router_058_src_valid),                                                  //          .valid
		.src_data           (id_router_058_src_data),                                                   //          .data
		.src_channel        (id_router_058_src_channel),                                                //          .channel
		.src_startofpacket  (id_router_058_src_startofpacket),                                          //          .startofpacket
		.src_endofpacket    (id_router_058_src_endofpacket)                                             //          .endofpacket
	);

	NIOS_SYSTEMV3_id_router_003 id_router_059 (
		.sink_ready         (ch2_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ch2_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ch2_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ch2_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ch2_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                  //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                       // clk_reset.reset
		.src_ready          (id_router_059_src_ready),                                                  //       src.ready
		.src_valid          (id_router_059_src_valid),                                                  //          .valid
		.src_data           (id_router_059_src_data),                                                   //          .data
		.src_channel        (id_router_059_src_channel),                                                //          .channel
		.src_startofpacket  (id_router_059_src_startofpacket),                                          //          .startofpacket
		.src_endofpacket    (id_router_059_src_endofpacket)                                             //          .endofpacket
	);

	NIOS_SYSTEMV3_id_router_003 id_router_060 (
		.sink_ready         (ch2_yn2_l_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ch2_yn2_l_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ch2_yn2_l_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ch2_yn2_l_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ch2_yn2_l_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                 //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                      // clk_reset.reset
		.src_ready          (id_router_060_src_ready),                                                 //       src.ready
		.src_valid          (id_router_060_src_valid),                                                 //          .valid
		.src_data           (id_router_060_src_data),                                                  //          .data
		.src_channel        (id_router_060_src_channel),                                               //          .channel
		.src_startofpacket  (id_router_060_src_startofpacket),                                         //          .startofpacket
		.src_endofpacket    (id_router_060_src_endofpacket)                                            //          .endofpacket
	);

	NIOS_SYSTEMV3_id_router_003 id_router_061 (
		.sink_ready         (ch2_yn3_u_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ch2_yn3_u_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ch2_yn3_u_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ch2_yn3_u_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ch2_yn3_u_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                 //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                      // clk_reset.reset
		.src_ready          (id_router_061_src_ready),                                                 //       src.ready
		.src_valid          (id_router_061_src_valid),                                                 //          .valid
		.src_data           (id_router_061_src_data),                                                  //          .data
		.src_channel        (id_router_061_src_channel),                                               //          .channel
		.src_startofpacket  (id_router_061_src_startofpacket),                                         //          .startofpacket
		.src_endofpacket    (id_router_061_src_endofpacket)                                            //          .endofpacket
	);

	NIOS_SYSTEMV3_id_router_003 id_router_062 (
		.sink_ready         (ch2_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ch2_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ch2_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ch2_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ch2_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                  //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                       // clk_reset.reset
		.src_ready          (id_router_062_src_ready),                                                  //       src.ready
		.src_valid          (id_router_062_src_valid),                                                  //          .valid
		.src_data           (id_router_062_src_data),                                                   //          .data
		.src_channel        (id_router_062_src_channel),                                                //          .channel
		.src_startofpacket  (id_router_062_src_startofpacket),                                          //          .startofpacket
		.src_endofpacket    (id_router_062_src_endofpacket)                                             //          .endofpacket
	);

	NIOS_SYSTEMV3_id_router_003 id_router_063 (
		.sink_ready         (ch2_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ch2_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ch2_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ch2_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ch2_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                  //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                       // clk_reset.reset
		.src_ready          (id_router_063_src_ready),                                                  //       src.ready
		.src_valid          (id_router_063_src_valid),                                                  //          .valid
		.src_data           (id_router_063_src_data),                                                   //          .data
		.src_channel        (id_router_063_src_channel),                                                //          .channel
		.src_startofpacket  (id_router_063_src_startofpacket),                                          //          .startofpacket
		.src_endofpacket    (id_router_063_src_endofpacket)                                             //          .endofpacket
	);

	NIOS_SYSTEMV3_id_router_003 id_router_064 (
		.sink_ready         (ch2_yn3_l_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ch2_yn3_l_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ch2_yn3_l_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ch2_yn3_l_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ch2_yn3_l_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                 //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                      // clk_reset.reset
		.src_ready          (id_router_064_src_ready),                                                 //       src.ready
		.src_valid          (id_router_064_src_valid),                                                 //          .valid
		.src_data           (id_router_064_src_data),                                                  //          .data
		.src_channel        (id_router_064_src_channel),                                               //          .channel
		.src_startofpacket  (id_router_064_src_startofpacket),                                         //          .startofpacket
		.src_endofpacket    (id_router_064_src_endofpacket)                                            //          .endofpacket
	);

	NIOS_SYSTEMV3_id_router_003 id_router_065 (
		.sink_ready         (ch3_timer_rst_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ch3_timer_rst_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ch3_timer_rst_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ch3_timer_rst_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ch3_timer_rst_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                     //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                          // clk_reset.reset
		.src_ready          (id_router_065_src_ready),                                                     //       src.ready
		.src_valid          (id_router_065_src_valid),                                                     //          .valid
		.src_data           (id_router_065_src_data),                                                      //          .data
		.src_channel        (id_router_065_src_channel),                                                   //          .channel
		.src_startofpacket  (id_router_065_src_startofpacket),                                             //          .startofpacket
		.src_endofpacket    (id_router_065_src_endofpacket)                                                //          .endofpacket
	);

	NIOS_SYSTEMV3_id_router_003 id_router_066 (
		.sink_ready         (ch3_thresh_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ch3_thresh_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ch3_thresh_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ch3_thresh_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ch3_thresh_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                  //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                       // clk_reset.reset
		.src_ready          (id_router_066_src_ready),                                                  //       src.ready
		.src_valid          (id_router_066_src_valid),                                                  //          .valid
		.src_data           (id_router_066_src_data),                                                   //          .data
		.src_channel        (id_router_066_src_channel),                                                //          .channel
		.src_startofpacket  (id_router_066_src_startofpacket),                                          //          .startofpacket
		.src_endofpacket    (id_router_066_src_endofpacket)                                             //          .endofpacket
	);

	NIOS_SYSTEMV3_id_router_003 id_router_067 (
		.sink_ready         (ch3_rd_peak_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ch3_rd_peak_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ch3_rd_peak_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ch3_rd_peak_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ch3_rd_peak_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                   //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                        // clk_reset.reset
		.src_ready          (id_router_067_src_ready),                                                   //       src.ready
		.src_valid          (id_router_067_src_valid),                                                   //          .valid
		.src_data           (id_router_067_src_data),                                                    //          .data
		.src_channel        (id_router_067_src_channel),                                                 //          .channel
		.src_startofpacket  (id_router_067_src_startofpacket),                                           //          .startofpacket
		.src_endofpacket    (id_router_067_src_endofpacket)                                              //          .endofpacket
	);

	NIOS_SYSTEMV3_id_router_003 id_router_068 (
		.sink_ready         (ch3_peak_found_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ch3_peak_found_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ch3_peak_found_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ch3_peak_found_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ch3_peak_found_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                      //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                           // clk_reset.reset
		.src_ready          (id_router_068_src_ready),                                                      //       src.ready
		.src_valid          (id_router_068_src_valid),                                                      //          .valid
		.src_data           (id_router_068_src_data),                                                       //          .data
		.src_channel        (id_router_068_src_channel),                                                    //          .channel
		.src_startofpacket  (id_router_068_src_startofpacket),                                              //          .startofpacket
		.src_endofpacket    (id_router_068_src_endofpacket)                                                 //          .endofpacket
	);

	NIOS_SYSTEMV3_id_router_003 id_router_069 (
		.sink_ready         (ch3_yn1_u_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ch3_yn1_u_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ch3_yn1_u_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ch3_yn1_u_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ch3_yn1_u_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                 //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                      // clk_reset.reset
		.src_ready          (id_router_069_src_ready),                                                 //       src.ready
		.src_valid          (id_router_069_src_valid),                                                 //          .valid
		.src_data           (id_router_069_src_data),                                                  //          .data
		.src_channel        (id_router_069_src_channel),                                               //          .channel
		.src_startofpacket  (id_router_069_src_startofpacket),                                         //          .startofpacket
		.src_endofpacket    (id_router_069_src_endofpacket)                                            //          .endofpacket
	);

	NIOS_SYSTEMV3_id_router_003 id_router_070 (
		.sink_ready         (ch3_time_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ch3_time_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ch3_time_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ch3_time_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ch3_time_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                     // clk_reset.reset
		.src_ready          (id_router_070_src_ready),                                                //       src.ready
		.src_valid          (id_router_070_src_valid),                                                //          .valid
		.src_data           (id_router_070_src_data),                                                 //          .data
		.src_channel        (id_router_070_src_channel),                                              //          .channel
		.src_startofpacket  (id_router_070_src_startofpacket),                                        //          .startofpacket
		.src_endofpacket    (id_router_070_src_endofpacket)                                           //          .endofpacket
	);

	NIOS_SYSTEMV3_id_router_003 id_router_071 (
		.sink_ready         (ch3_yn3_l_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ch3_yn3_l_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ch3_yn3_l_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ch3_yn3_l_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ch3_yn3_l_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                 //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                      // clk_reset.reset
		.src_ready          (id_router_071_src_ready),                                                 //       src.ready
		.src_valid          (id_router_071_src_valid),                                                 //          .valid
		.src_data           (id_router_071_src_data),                                                  //          .data
		.src_channel        (id_router_071_src_channel),                                               //          .channel
		.src_startofpacket  (id_router_071_src_startofpacket),                                         //          .startofpacket
		.src_endofpacket    (id_router_071_src_endofpacket)                                            //          .endofpacket
	);

	NIOS_SYSTEMV3_id_router_003 id_router_072 (
		.sink_ready         (ch3_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ch3_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ch3_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ch3_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ch3_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                  //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                       // clk_reset.reset
		.src_ready          (id_router_072_src_ready),                                                  //       src.ready
		.src_valid          (id_router_072_src_valid),                                                  //          .valid
		.src_data           (id_router_072_src_data),                                                   //          .data
		.src_channel        (id_router_072_src_channel),                                                //          .channel
		.src_startofpacket  (id_router_072_src_startofpacket),                                          //          .startofpacket
		.src_endofpacket    (id_router_072_src_endofpacket)                                             //          .endofpacket
	);

	NIOS_SYSTEMV3_id_router_003 id_router_073 (
		.sink_ready         (ch3_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ch3_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ch3_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ch3_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ch3_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                  //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                       // clk_reset.reset
		.src_ready          (id_router_073_src_ready),                                                  //       src.ready
		.src_valid          (id_router_073_src_valid),                                                  //          .valid
		.src_data           (id_router_073_src_data),                                                   //          .data
		.src_channel        (id_router_073_src_channel),                                                //          .channel
		.src_startofpacket  (id_router_073_src_startofpacket),                                          //          .startofpacket
		.src_endofpacket    (id_router_073_src_endofpacket)                                             //          .endofpacket
	);

	NIOS_SYSTEMV3_id_router_003 id_router_074 (
		.sink_ready         (ch3_yn3_u_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ch3_yn3_u_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ch3_yn3_u_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ch3_yn3_u_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ch3_yn3_u_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                 //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                      // clk_reset.reset
		.src_ready          (id_router_074_src_ready),                                                 //       src.ready
		.src_valid          (id_router_074_src_valid),                                                 //          .valid
		.src_data           (id_router_074_src_data),                                                  //          .data
		.src_channel        (id_router_074_src_channel),                                               //          .channel
		.src_startofpacket  (id_router_074_src_startofpacket),                                         //          .startofpacket
		.src_endofpacket    (id_router_074_src_endofpacket)                                            //          .endofpacket
	);

	NIOS_SYSTEMV3_id_router_003 id_router_075 (
		.sink_ready         (ch3_yn2_l_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ch3_yn2_l_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ch3_yn2_l_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ch3_yn2_l_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ch3_yn2_l_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                 //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                      // clk_reset.reset
		.src_ready          (id_router_075_src_ready),                                                 //       src.ready
		.src_valid          (id_router_075_src_valid),                                                 //          .valid
		.src_data           (id_router_075_src_data),                                                  //          .data
		.src_channel        (id_router_075_src_channel),                                               //          .channel
		.src_startofpacket  (id_router_075_src_startofpacket),                                         //          .startofpacket
		.src_endofpacket    (id_router_075_src_endofpacket)                                            //          .endofpacket
	);

	NIOS_SYSTEMV3_id_router_003 id_router_076 (
		.sink_ready         (ch3_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ch3_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ch3_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ch3_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ch3_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                  //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                       // clk_reset.reset
		.src_ready          (id_router_076_src_ready),                                                  //       src.ready
		.src_valid          (id_router_076_src_valid),                                                  //          .valid
		.src_data           (id_router_076_src_data),                                                   //          .data
		.src_channel        (id_router_076_src_channel),                                                //          .channel
		.src_startofpacket  (id_router_076_src_startofpacket),                                          //          .startofpacket
		.src_endofpacket    (id_router_076_src_endofpacket)                                             //          .endofpacket
	);

	NIOS_SYSTEMV3_id_router_003 id_router_077 (
		.sink_ready         (ch3_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ch3_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ch3_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ch3_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ch3_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                  //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                       // clk_reset.reset
		.src_ready          (id_router_077_src_ready),                                                  //       src.ready
		.src_valid          (id_router_077_src_valid),                                                  //          .valid
		.src_data           (id_router_077_src_data),                                                   //          .data
		.src_channel        (id_router_077_src_channel),                                                //          .channel
		.src_startofpacket  (id_router_077_src_startofpacket),                                          //          .startofpacket
		.src_endofpacket    (id_router_077_src_endofpacket)                                             //          .endofpacket
	);

	NIOS_SYSTEMV3_id_router_003 id_router_078 (
		.sink_ready         (ch3_yn2_u_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ch3_yn2_u_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ch3_yn2_u_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ch3_yn2_u_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ch3_yn2_u_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                 //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                      // clk_reset.reset
		.src_ready          (id_router_078_src_ready),                                                 //       src.ready
		.src_valid          (id_router_078_src_valid),                                                 //          .valid
		.src_data           (id_router_078_src_data),                                                  //          .data
		.src_channel        (id_router_078_src_channel),                                               //          .channel
		.src_startofpacket  (id_router_078_src_startofpacket),                                         //          .startofpacket
		.src_endofpacket    (id_router_078_src_endofpacket)                                            //          .endofpacket
	);

	NIOS_SYSTEMV3_id_router_003 id_router_079 (
		.sink_ready         (ch3_yn1_l_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ch3_yn1_l_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ch3_yn1_l_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ch3_yn1_l_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ch3_yn1_l_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                 //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                      // clk_reset.reset
		.src_ready          (id_router_079_src_ready),                                                 //       src.ready
		.src_valid          (id_router_079_src_valid),                                                 //          .valid
		.src_data           (id_router_079_src_data),                                                  //          .data
		.src_channel        (id_router_079_src_channel),                                               //          .channel
		.src_startofpacket  (id_router_079_src_startofpacket),                                         //          .startofpacket
		.src_endofpacket    (id_router_079_src_endofpacket)                                            //          .endofpacket
	);

	NIOS_SYSTEMV3_id_router_003 id_router_080 (
		.sink_ready         (ch3_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ch3_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ch3_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ch3_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ch3_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                  //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                       // clk_reset.reset
		.src_ready          (id_router_080_src_ready),                                                  //       src.ready
		.src_valid          (id_router_080_src_valid),                                                  //          .valid
		.src_data           (id_router_080_src_data),                                                   //          .data
		.src_channel        (id_router_080_src_channel),                                                //          .channel
		.src_startofpacket  (id_router_080_src_startofpacket),                                          //          .startofpacket
		.src_endofpacket    (id_router_080_src_endofpacket)                                             //          .endofpacket
	);

	NIOS_SYSTEMV3_id_router_003 id_router_081 (
		.sink_ready         (ch3_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ch3_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ch3_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ch3_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ch3_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                  //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                       // clk_reset.reset
		.src_ready          (id_router_081_src_ready),                                                  //       src.ready
		.src_valid          (id_router_081_src_valid),                                                  //          .valid
		.src_data           (id_router_081_src_data),                                                   //          .data
		.src_channel        (id_router_081_src_channel),                                                //          .channel
		.src_startofpacket  (id_router_081_src_startofpacket),                                          //          .startofpacket
		.src_endofpacket    (id_router_081_src_endofpacket)                                             //          .endofpacket
	);

	NIOS_SYSTEMV3_id_router_003 id_router_082 (
		.sink_ready         (ch4_timer_rst_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ch4_timer_rst_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ch4_timer_rst_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ch4_timer_rst_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ch4_timer_rst_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                     //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                          // clk_reset.reset
		.src_ready          (id_router_082_src_ready),                                                     //       src.ready
		.src_valid          (id_router_082_src_valid),                                                     //          .valid
		.src_data           (id_router_082_src_data),                                                      //          .data
		.src_channel        (id_router_082_src_channel),                                                   //          .channel
		.src_startofpacket  (id_router_082_src_startofpacket),                                             //          .startofpacket
		.src_endofpacket    (id_router_082_src_endofpacket)                                                //          .endofpacket
	);

	NIOS_SYSTEMV3_id_router_003 id_router_083 (
		.sink_ready         (ch4_thresh_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ch4_thresh_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ch4_thresh_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ch4_thresh_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ch4_thresh_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                  //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                       // clk_reset.reset
		.src_ready          (id_router_083_src_ready),                                                  //       src.ready
		.src_valid          (id_router_083_src_valid),                                                  //          .valid
		.src_data           (id_router_083_src_data),                                                   //          .data
		.src_channel        (id_router_083_src_channel),                                                //          .channel
		.src_startofpacket  (id_router_083_src_startofpacket),                                          //          .startofpacket
		.src_endofpacket    (id_router_083_src_endofpacket)                                             //          .endofpacket
	);

	NIOS_SYSTEMV3_id_router_003 id_router_084 (
		.sink_ready         (ch4_rd_peak_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ch4_rd_peak_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ch4_rd_peak_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ch4_rd_peak_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ch4_rd_peak_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                   //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                        // clk_reset.reset
		.src_ready          (id_router_084_src_ready),                                                   //       src.ready
		.src_valid          (id_router_084_src_valid),                                                   //          .valid
		.src_data           (id_router_084_src_data),                                                    //          .data
		.src_channel        (id_router_084_src_channel),                                                 //          .channel
		.src_startofpacket  (id_router_084_src_startofpacket),                                           //          .startofpacket
		.src_endofpacket    (id_router_084_src_endofpacket)                                              //          .endofpacket
	);

	NIOS_SYSTEMV3_id_router_003 id_router_085 (
		.sink_ready         (ch4_peak_found_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ch4_peak_found_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ch4_peak_found_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ch4_peak_found_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ch4_peak_found_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                      //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                           // clk_reset.reset
		.src_ready          (id_router_085_src_ready),                                                      //       src.ready
		.src_valid          (id_router_085_src_valid),                                                      //          .valid
		.src_data           (id_router_085_src_data),                                                       //          .data
		.src_channel        (id_router_085_src_channel),                                                    //          .channel
		.src_startofpacket  (id_router_085_src_startofpacket),                                              //          .startofpacket
		.src_endofpacket    (id_router_085_src_endofpacket)                                                 //          .endofpacket
	);

	NIOS_SYSTEMV3_id_router_003 id_router_086 (
		.sink_ready         (ch4_time_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ch4_time_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ch4_time_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ch4_time_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ch4_time_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                     // clk_reset.reset
		.src_ready          (id_router_086_src_ready),                                                //       src.ready
		.src_valid          (id_router_086_src_valid),                                                //          .valid
		.src_data           (id_router_086_src_data),                                                 //          .data
		.src_channel        (id_router_086_src_channel),                                              //          .channel
		.src_startofpacket  (id_router_086_src_startofpacket),                                        //          .startofpacket
		.src_endofpacket    (id_router_086_src_endofpacket)                                           //          .endofpacket
	);

	NIOS_SYSTEMV3_id_router_003 id_router_087 (
		.sink_ready         (ch4_yn1_u_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ch4_yn1_u_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ch4_yn1_u_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ch4_yn1_u_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ch4_yn1_u_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                 //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                      // clk_reset.reset
		.src_ready          (id_router_087_src_ready),                                                 //       src.ready
		.src_valid          (id_router_087_src_valid),                                                 //          .valid
		.src_data           (id_router_087_src_data),                                                  //          .data
		.src_channel        (id_router_087_src_channel),                                               //          .channel
		.src_startofpacket  (id_router_087_src_startofpacket),                                         //          .startofpacket
		.src_endofpacket    (id_router_087_src_endofpacket)                                            //          .endofpacket
	);

	NIOS_SYSTEMV3_id_router_003 id_router_088 (
		.sink_ready         (ch4_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ch4_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ch4_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ch4_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ch4_yn1_mu_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                  //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                       // clk_reset.reset
		.src_ready          (id_router_088_src_ready),                                                  //       src.ready
		.src_valid          (id_router_088_src_valid),                                                  //          .valid
		.src_data           (id_router_088_src_data),                                                   //          .data
		.src_channel        (id_router_088_src_channel),                                                //          .channel
		.src_startofpacket  (id_router_088_src_startofpacket),                                          //          .startofpacket
		.src_endofpacket    (id_router_088_src_endofpacket)                                             //          .endofpacket
	);

	NIOS_SYSTEMV3_id_router_003 id_router_089 (
		.sink_ready         (ch4_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ch4_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ch4_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ch4_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ch4_yn1_ml_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                  //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                       // clk_reset.reset
		.src_ready          (id_router_089_src_ready),                                                  //       src.ready
		.src_valid          (id_router_089_src_valid),                                                  //          .valid
		.src_data           (id_router_089_src_data),                                                   //          .data
		.src_channel        (id_router_089_src_channel),                                                //          .channel
		.src_startofpacket  (id_router_089_src_startofpacket),                                          //          .startofpacket
		.src_endofpacket    (id_router_089_src_endofpacket)                                             //          .endofpacket
	);

	NIOS_SYSTEMV3_id_router_003 id_router_090 (
		.sink_ready         (ch4_yn1_l_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ch4_yn1_l_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ch4_yn1_l_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ch4_yn1_l_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ch4_yn1_l_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                 //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                      // clk_reset.reset
		.src_ready          (id_router_090_src_ready),                                                 //       src.ready
		.src_valid          (id_router_090_src_valid),                                                 //          .valid
		.src_data           (id_router_090_src_data),                                                  //          .data
		.src_channel        (id_router_090_src_channel),                                               //          .channel
		.src_startofpacket  (id_router_090_src_startofpacket),                                         //          .startofpacket
		.src_endofpacket    (id_router_090_src_endofpacket)                                            //          .endofpacket
	);

	NIOS_SYSTEMV3_id_router_003 id_router_091 (
		.sink_ready         (ch4_yn2_u_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ch4_yn2_u_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ch4_yn2_u_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ch4_yn2_u_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ch4_yn2_u_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                 //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                      // clk_reset.reset
		.src_ready          (id_router_091_src_ready),                                                 //       src.ready
		.src_valid          (id_router_091_src_valid),                                                 //          .valid
		.src_data           (id_router_091_src_data),                                                  //          .data
		.src_channel        (id_router_091_src_channel),                                               //          .channel
		.src_startofpacket  (id_router_091_src_startofpacket),                                         //          .startofpacket
		.src_endofpacket    (id_router_091_src_endofpacket)                                            //          .endofpacket
	);

	NIOS_SYSTEMV3_id_router_003 id_router_092 (
		.sink_ready         (ch4_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ch4_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ch4_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ch4_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ch4_yn2_mu_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                  //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                       // clk_reset.reset
		.src_ready          (id_router_092_src_ready),                                                  //       src.ready
		.src_valid          (id_router_092_src_valid),                                                  //          .valid
		.src_data           (id_router_092_src_data),                                                   //          .data
		.src_channel        (id_router_092_src_channel),                                                //          .channel
		.src_startofpacket  (id_router_092_src_startofpacket),                                          //          .startofpacket
		.src_endofpacket    (id_router_092_src_endofpacket)                                             //          .endofpacket
	);

	NIOS_SYSTEMV3_id_router_003 id_router_093 (
		.sink_ready         (ch4_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ch4_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ch4_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ch4_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ch4_yn2_ml_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                  //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                       // clk_reset.reset
		.src_ready          (id_router_093_src_ready),                                                  //       src.ready
		.src_valid          (id_router_093_src_valid),                                                  //          .valid
		.src_data           (id_router_093_src_data),                                                   //          .data
		.src_channel        (id_router_093_src_channel),                                                //          .channel
		.src_startofpacket  (id_router_093_src_startofpacket),                                          //          .startofpacket
		.src_endofpacket    (id_router_093_src_endofpacket)                                             //          .endofpacket
	);

	NIOS_SYSTEMV3_id_router_003 id_router_094 (
		.sink_ready         (ch4_yn2_l_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ch4_yn2_l_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ch4_yn2_l_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ch4_yn2_l_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ch4_yn2_l_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                 //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                      // clk_reset.reset
		.src_ready          (id_router_094_src_ready),                                                 //       src.ready
		.src_valid          (id_router_094_src_valid),                                                 //          .valid
		.src_data           (id_router_094_src_data),                                                  //          .data
		.src_channel        (id_router_094_src_channel),                                               //          .channel
		.src_startofpacket  (id_router_094_src_startofpacket),                                         //          .startofpacket
		.src_endofpacket    (id_router_094_src_endofpacket)                                            //          .endofpacket
	);

	NIOS_SYSTEMV3_id_router_003 id_router_095 (
		.sink_ready         (ch4_yn3_u_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ch4_yn3_u_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ch4_yn3_u_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ch4_yn3_u_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ch4_yn3_u_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                 //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                      // clk_reset.reset
		.src_ready          (id_router_095_src_ready),                                                 //       src.ready
		.src_valid          (id_router_095_src_valid),                                                 //          .valid
		.src_data           (id_router_095_src_data),                                                  //          .data
		.src_channel        (id_router_095_src_channel),                                               //          .channel
		.src_startofpacket  (id_router_095_src_startofpacket),                                         //          .startofpacket
		.src_endofpacket    (id_router_095_src_endofpacket)                                            //          .endofpacket
	);

	NIOS_SYSTEMV3_id_router_003 id_router_096 (
		.sink_ready         (ch4_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ch4_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ch4_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ch4_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ch4_yn3_mu_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                  //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                       // clk_reset.reset
		.src_ready          (id_router_096_src_ready),                                                  //       src.ready
		.src_valid          (id_router_096_src_valid),                                                  //          .valid
		.src_data           (id_router_096_src_data),                                                   //          .data
		.src_channel        (id_router_096_src_channel),                                                //          .channel
		.src_startofpacket  (id_router_096_src_startofpacket),                                          //          .startofpacket
		.src_endofpacket    (id_router_096_src_endofpacket)                                             //          .endofpacket
	);

	NIOS_SYSTEMV3_id_router_003 id_router_097 (
		.sink_ready         (ch4_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ch4_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ch4_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ch4_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ch4_yn3_ml_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                  //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                       // clk_reset.reset
		.src_ready          (id_router_097_src_ready),                                                  //       src.ready
		.src_valid          (id_router_097_src_valid),                                                  //          .valid
		.src_data           (id_router_097_src_data),                                                   //          .data
		.src_channel        (id_router_097_src_channel),                                                //          .channel
		.src_startofpacket  (id_router_097_src_startofpacket),                                          //          .startofpacket
		.src_endofpacket    (id_router_097_src_endofpacket)                                             //          .endofpacket
	);

	NIOS_SYSTEMV3_id_router_003 id_router_098 (
		.sink_ready         (ch4_yn3_l_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ch4_yn3_l_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ch4_yn3_l_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ch4_yn3_l_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ch4_yn3_l_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                 //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                      // clk_reset.reset
		.src_ready          (id_router_098_src_ready),                                                 //       src.ready
		.src_valid          (id_router_098_src_valid),                                                 //          .valid
		.src_data           (id_router_098_src_data),                                                  //          .data
		.src_channel        (id_router_098_src_channel),                                               //          .channel
		.src_startofpacket  (id_router_098_src_startofpacket),                                         //          .startofpacket
		.src_endofpacket    (id_router_098_src_endofpacket)                                            //          .endofpacket
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (1),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2),
		.RESET_REQUEST_PRESENT   (0)
	) rst_controller (
		.reset_in0  (~reset_reset_n),                 // reset_in0.reset
		.clk        (clk_clk),                        //       clk.clk
		.reset_out  (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req  (),                               // (terminated)
		.reset_in1  (1'b0),                           // (terminated)
		.reset_in2  (1'b0),                           // (terminated)
		.reset_in3  (1'b0),                           // (terminated)
		.reset_in4  (1'b0),                           // (terminated)
		.reset_in5  (1'b0),                           // (terminated)
		.reset_in6  (1'b0),                           // (terminated)
		.reset_in7  (1'b0),                           // (terminated)
		.reset_in8  (1'b0),                           // (terminated)
		.reset_in9  (1'b0),                           // (terminated)
		.reset_in10 (1'b0),                           // (terminated)
		.reset_in11 (1'b0),                           // (terminated)
		.reset_in12 (1'b0),                           // (terminated)
		.reset_in13 (1'b0),                           // (terminated)
		.reset_in14 (1'b0),                           // (terminated)
		.reset_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (2),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2),
		.RESET_REQUEST_PRESENT   (1)
	) rst_controller_001 (
		.reset_in0  (nios_cpu_jtag_debug_module_reset_reset), // reset_in0.reset
		.reset_in1  (~reset_reset_n),                         // reset_in1.reset
		.clk        (clk_clk),                                //       clk.clk
		.reset_out  (rst_controller_001_reset_out_reset),     // reset_out.reset
		.reset_req  (rst_controller_001_reset_out_reset_req), //          .reset_req
		.reset_in2  (1'b0),                                   // (terminated)
		.reset_in3  (1'b0),                                   // (terminated)
		.reset_in4  (1'b0),                                   // (terminated)
		.reset_in5  (1'b0),                                   // (terminated)
		.reset_in6  (1'b0),                                   // (terminated)
		.reset_in7  (1'b0),                                   // (terminated)
		.reset_in8  (1'b0),                                   // (terminated)
		.reset_in9  (1'b0),                                   // (terminated)
		.reset_in10 (1'b0),                                   // (terminated)
		.reset_in11 (1'b0),                                   // (terminated)
		.reset_in12 (1'b0),                                   // (terminated)
		.reset_in13 (1'b0),                                   // (terminated)
		.reset_in14 (1'b0),                                   // (terminated)
		.reset_in15 (1'b0)                                    // (terminated)
	);

	NIOS_SYSTEMV3_cmd_xbar_demux cmd_xbar_demux (
		.clk                (clk_clk),                           //       clk.clk
		.reset              (rst_controller_reset_out_reset),    // clk_reset.reset
		.sink_ready         (addr_router_src_ready),             //      sink.ready
		.sink_channel       (addr_router_src_channel),           //          .channel
		.sink_data          (addr_router_src_data),              //          .data
		.sink_startofpacket (addr_router_src_startofpacket),     //          .startofpacket
		.sink_endofpacket   (addr_router_src_endofpacket),       //          .endofpacket
		.sink_valid         (addr_router_src_valid),             //          .valid
		.src0_ready         (cmd_xbar_demux_src0_ready),         //      src0.ready
		.src0_valid         (cmd_xbar_demux_src0_valid),         //          .valid
		.src0_data          (cmd_xbar_demux_src0_data),          //          .data
		.src0_channel       (cmd_xbar_demux_src0_channel),       //          .channel
		.src0_startofpacket (cmd_xbar_demux_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_src0_endofpacket),   //          .endofpacket
		.src1_ready         (cmd_xbar_demux_src1_ready),         //      src1.ready
		.src1_valid         (cmd_xbar_demux_src1_valid),         //          .valid
		.src1_data          (cmd_xbar_demux_src1_data),          //          .data
		.src1_channel       (cmd_xbar_demux_src1_channel),       //          .channel
		.src1_startofpacket (cmd_xbar_demux_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (cmd_xbar_demux_src1_endofpacket),   //          .endofpacket
		.src2_ready         (cmd_xbar_demux_src2_ready),         //      src2.ready
		.src2_valid         (cmd_xbar_demux_src2_valid),         //          .valid
		.src2_data          (cmd_xbar_demux_src2_data),          //          .data
		.src2_channel       (cmd_xbar_demux_src2_channel),       //          .channel
		.src2_startofpacket (cmd_xbar_demux_src2_startofpacket), //          .startofpacket
		.src2_endofpacket   (cmd_xbar_demux_src2_endofpacket)    //          .endofpacket
	);

	NIOS_SYSTEMV3_cmd_xbar_demux_001 cmd_xbar_demux_001 (
		.clk                 (clk_clk),                                //       clk.clk
		.reset               (rst_controller_reset_out_reset),         // clk_reset.reset
		.sink_ready          (addr_router_001_src_ready),              //      sink.ready
		.sink_channel        (addr_router_001_src_channel),            //          .channel
		.sink_data           (addr_router_001_src_data),               //          .data
		.sink_startofpacket  (addr_router_001_src_startofpacket),      //          .startofpacket
		.sink_endofpacket    (addr_router_001_src_endofpacket),        //          .endofpacket
		.sink_valid          (addr_router_001_src_valid),              //          .valid
		.src0_ready          (cmd_xbar_demux_001_src0_ready),          //      src0.ready
		.src0_valid          (cmd_xbar_demux_001_src0_valid),          //          .valid
		.src0_data           (cmd_xbar_demux_001_src0_data),           //          .data
		.src0_channel        (cmd_xbar_demux_001_src0_channel),        //          .channel
		.src0_startofpacket  (cmd_xbar_demux_001_src0_startofpacket),  //          .startofpacket
		.src0_endofpacket    (cmd_xbar_demux_001_src0_endofpacket),    //          .endofpacket
		.src1_ready          (cmd_xbar_demux_001_src1_ready),          //      src1.ready
		.src1_valid          (cmd_xbar_demux_001_src1_valid),          //          .valid
		.src1_data           (cmd_xbar_demux_001_src1_data),           //          .data
		.src1_channel        (cmd_xbar_demux_001_src1_channel),        //          .channel
		.src1_startofpacket  (cmd_xbar_demux_001_src1_startofpacket),  //          .startofpacket
		.src1_endofpacket    (cmd_xbar_demux_001_src1_endofpacket),    //          .endofpacket
		.src2_ready          (cmd_xbar_demux_001_src2_ready),          //      src2.ready
		.src2_valid          (cmd_xbar_demux_001_src2_valid),          //          .valid
		.src2_data           (cmd_xbar_demux_001_src2_data),           //          .data
		.src2_channel        (cmd_xbar_demux_001_src2_channel),        //          .channel
		.src2_startofpacket  (cmd_xbar_demux_001_src2_startofpacket),  //          .startofpacket
		.src2_endofpacket    (cmd_xbar_demux_001_src2_endofpacket),    //          .endofpacket
		.src3_ready          (cmd_xbar_demux_001_src3_ready),          //      src3.ready
		.src3_valid          (cmd_xbar_demux_001_src3_valid),          //          .valid
		.src3_data           (cmd_xbar_demux_001_src3_data),           //          .data
		.src3_channel        (cmd_xbar_demux_001_src3_channel),        //          .channel
		.src3_startofpacket  (cmd_xbar_demux_001_src3_startofpacket),  //          .startofpacket
		.src3_endofpacket    (cmd_xbar_demux_001_src3_endofpacket),    //          .endofpacket
		.src4_ready          (cmd_xbar_demux_001_src4_ready),          //      src4.ready
		.src4_valid          (cmd_xbar_demux_001_src4_valid),          //          .valid
		.src4_data           (cmd_xbar_demux_001_src4_data),           //          .data
		.src4_channel        (cmd_xbar_demux_001_src4_channel),        //          .channel
		.src4_startofpacket  (cmd_xbar_demux_001_src4_startofpacket),  //          .startofpacket
		.src4_endofpacket    (cmd_xbar_demux_001_src4_endofpacket),    //          .endofpacket
		.src5_ready          (cmd_xbar_demux_001_src5_ready),          //      src5.ready
		.src5_valid          (cmd_xbar_demux_001_src5_valid),          //          .valid
		.src5_data           (cmd_xbar_demux_001_src5_data),           //          .data
		.src5_channel        (cmd_xbar_demux_001_src5_channel),        //          .channel
		.src5_startofpacket  (cmd_xbar_demux_001_src5_startofpacket),  //          .startofpacket
		.src5_endofpacket    (cmd_xbar_demux_001_src5_endofpacket),    //          .endofpacket
		.src6_ready          (cmd_xbar_demux_001_src6_ready),          //      src6.ready
		.src6_valid          (cmd_xbar_demux_001_src6_valid),          //          .valid
		.src6_data           (cmd_xbar_demux_001_src6_data),           //          .data
		.src6_channel        (cmd_xbar_demux_001_src6_channel),        //          .channel
		.src6_startofpacket  (cmd_xbar_demux_001_src6_startofpacket),  //          .startofpacket
		.src6_endofpacket    (cmd_xbar_demux_001_src6_endofpacket),    //          .endofpacket
		.src7_ready          (cmd_xbar_demux_001_src7_ready),          //      src7.ready
		.src7_valid          (cmd_xbar_demux_001_src7_valid),          //          .valid
		.src7_data           (cmd_xbar_demux_001_src7_data),           //          .data
		.src7_channel        (cmd_xbar_demux_001_src7_channel),        //          .channel
		.src7_startofpacket  (cmd_xbar_demux_001_src7_startofpacket),  //          .startofpacket
		.src7_endofpacket    (cmd_xbar_demux_001_src7_endofpacket),    //          .endofpacket
		.src8_ready          (cmd_xbar_demux_001_src8_ready),          //      src8.ready
		.src8_valid          (cmd_xbar_demux_001_src8_valid),          //          .valid
		.src8_data           (cmd_xbar_demux_001_src8_data),           //          .data
		.src8_channel        (cmd_xbar_demux_001_src8_channel),        //          .channel
		.src8_startofpacket  (cmd_xbar_demux_001_src8_startofpacket),  //          .startofpacket
		.src8_endofpacket    (cmd_xbar_demux_001_src8_endofpacket),    //          .endofpacket
		.src9_ready          (cmd_xbar_demux_001_src9_ready),          //      src9.ready
		.src9_valid          (cmd_xbar_demux_001_src9_valid),          //          .valid
		.src9_data           (cmd_xbar_demux_001_src9_data),           //          .data
		.src9_channel        (cmd_xbar_demux_001_src9_channel),        //          .channel
		.src9_startofpacket  (cmd_xbar_demux_001_src9_startofpacket),  //          .startofpacket
		.src9_endofpacket    (cmd_xbar_demux_001_src9_endofpacket),    //          .endofpacket
		.src10_ready         (cmd_xbar_demux_001_src10_ready),         //     src10.ready
		.src10_valid         (cmd_xbar_demux_001_src10_valid),         //          .valid
		.src10_data          (cmd_xbar_demux_001_src10_data),          //          .data
		.src10_channel       (cmd_xbar_demux_001_src10_channel),       //          .channel
		.src10_startofpacket (cmd_xbar_demux_001_src10_startofpacket), //          .startofpacket
		.src10_endofpacket   (cmd_xbar_demux_001_src10_endofpacket),   //          .endofpacket
		.src11_ready         (cmd_xbar_demux_001_src11_ready),         //     src11.ready
		.src11_valid         (cmd_xbar_demux_001_src11_valid),         //          .valid
		.src11_data          (cmd_xbar_demux_001_src11_data),          //          .data
		.src11_channel       (cmd_xbar_demux_001_src11_channel),       //          .channel
		.src11_startofpacket (cmd_xbar_demux_001_src11_startofpacket), //          .startofpacket
		.src11_endofpacket   (cmd_xbar_demux_001_src11_endofpacket),   //          .endofpacket
		.src12_ready         (cmd_xbar_demux_001_src12_ready),         //     src12.ready
		.src12_valid         (cmd_xbar_demux_001_src12_valid),         //          .valid
		.src12_data          (cmd_xbar_demux_001_src12_data),          //          .data
		.src12_channel       (cmd_xbar_demux_001_src12_channel),       //          .channel
		.src12_startofpacket (cmd_xbar_demux_001_src12_startofpacket), //          .startofpacket
		.src12_endofpacket   (cmd_xbar_demux_001_src12_endofpacket),   //          .endofpacket
		.src13_ready         (cmd_xbar_demux_001_src13_ready),         //     src13.ready
		.src13_valid         (cmd_xbar_demux_001_src13_valid),         //          .valid
		.src13_data          (cmd_xbar_demux_001_src13_data),          //          .data
		.src13_channel       (cmd_xbar_demux_001_src13_channel),       //          .channel
		.src13_startofpacket (cmd_xbar_demux_001_src13_startofpacket), //          .startofpacket
		.src13_endofpacket   (cmd_xbar_demux_001_src13_endofpacket),   //          .endofpacket
		.src14_ready         (cmd_xbar_demux_001_src14_ready),         //     src14.ready
		.src14_valid         (cmd_xbar_demux_001_src14_valid),         //          .valid
		.src14_data          (cmd_xbar_demux_001_src14_data),          //          .data
		.src14_channel       (cmd_xbar_demux_001_src14_channel),       //          .channel
		.src14_startofpacket (cmd_xbar_demux_001_src14_startofpacket), //          .startofpacket
		.src14_endofpacket   (cmd_xbar_demux_001_src14_endofpacket),   //          .endofpacket
		.src15_ready         (cmd_xbar_demux_001_src15_ready),         //     src15.ready
		.src15_valid         (cmd_xbar_demux_001_src15_valid),         //          .valid
		.src15_data          (cmd_xbar_demux_001_src15_data),          //          .data
		.src15_channel       (cmd_xbar_demux_001_src15_channel),       //          .channel
		.src15_startofpacket (cmd_xbar_demux_001_src15_startofpacket), //          .startofpacket
		.src15_endofpacket   (cmd_xbar_demux_001_src15_endofpacket),   //          .endofpacket
		.src16_ready         (cmd_xbar_demux_001_src16_ready),         //     src16.ready
		.src16_valid         (cmd_xbar_demux_001_src16_valid),         //          .valid
		.src16_data          (cmd_xbar_demux_001_src16_data),          //          .data
		.src16_channel       (cmd_xbar_demux_001_src16_channel),       //          .channel
		.src16_startofpacket (cmd_xbar_demux_001_src16_startofpacket), //          .startofpacket
		.src16_endofpacket   (cmd_xbar_demux_001_src16_endofpacket),   //          .endofpacket
		.src17_ready         (cmd_xbar_demux_001_src17_ready),         //     src17.ready
		.src17_valid         (cmd_xbar_demux_001_src17_valid),         //          .valid
		.src17_data          (cmd_xbar_demux_001_src17_data),          //          .data
		.src17_channel       (cmd_xbar_demux_001_src17_channel),       //          .channel
		.src17_startofpacket (cmd_xbar_demux_001_src17_startofpacket), //          .startofpacket
		.src17_endofpacket   (cmd_xbar_demux_001_src17_endofpacket),   //          .endofpacket
		.src18_ready         (cmd_xbar_demux_001_src18_ready),         //     src18.ready
		.src18_valid         (cmd_xbar_demux_001_src18_valid),         //          .valid
		.src18_data          (cmd_xbar_demux_001_src18_data),          //          .data
		.src18_channel       (cmd_xbar_demux_001_src18_channel),       //          .channel
		.src18_startofpacket (cmd_xbar_demux_001_src18_startofpacket), //          .startofpacket
		.src18_endofpacket   (cmd_xbar_demux_001_src18_endofpacket),   //          .endofpacket
		.src19_ready         (cmd_xbar_demux_001_src19_ready),         //     src19.ready
		.src19_valid         (cmd_xbar_demux_001_src19_valid),         //          .valid
		.src19_data          (cmd_xbar_demux_001_src19_data),          //          .data
		.src19_channel       (cmd_xbar_demux_001_src19_channel),       //          .channel
		.src19_startofpacket (cmd_xbar_demux_001_src19_startofpacket), //          .startofpacket
		.src19_endofpacket   (cmd_xbar_demux_001_src19_endofpacket),   //          .endofpacket
		.src20_ready         (cmd_xbar_demux_001_src20_ready),         //     src20.ready
		.src20_valid         (cmd_xbar_demux_001_src20_valid),         //          .valid
		.src20_data          (cmd_xbar_demux_001_src20_data),          //          .data
		.src20_channel       (cmd_xbar_demux_001_src20_channel),       //          .channel
		.src20_startofpacket (cmd_xbar_demux_001_src20_startofpacket), //          .startofpacket
		.src20_endofpacket   (cmd_xbar_demux_001_src20_endofpacket),   //          .endofpacket
		.src21_ready         (cmd_xbar_demux_001_src21_ready),         //     src21.ready
		.src21_valid         (cmd_xbar_demux_001_src21_valid),         //          .valid
		.src21_data          (cmd_xbar_demux_001_src21_data),          //          .data
		.src21_channel       (cmd_xbar_demux_001_src21_channel),       //          .channel
		.src21_startofpacket (cmd_xbar_demux_001_src21_startofpacket), //          .startofpacket
		.src21_endofpacket   (cmd_xbar_demux_001_src21_endofpacket),   //          .endofpacket
		.src22_ready         (cmd_xbar_demux_001_src22_ready),         //     src22.ready
		.src22_valid         (cmd_xbar_demux_001_src22_valid),         //          .valid
		.src22_data          (cmd_xbar_demux_001_src22_data),          //          .data
		.src22_channel       (cmd_xbar_demux_001_src22_channel),       //          .channel
		.src22_startofpacket (cmd_xbar_demux_001_src22_startofpacket), //          .startofpacket
		.src22_endofpacket   (cmd_xbar_demux_001_src22_endofpacket),   //          .endofpacket
		.src23_ready         (cmd_xbar_demux_001_src23_ready),         //     src23.ready
		.src23_valid         (cmd_xbar_demux_001_src23_valid),         //          .valid
		.src23_data          (cmd_xbar_demux_001_src23_data),          //          .data
		.src23_channel       (cmd_xbar_demux_001_src23_channel),       //          .channel
		.src23_startofpacket (cmd_xbar_demux_001_src23_startofpacket), //          .startofpacket
		.src23_endofpacket   (cmd_xbar_demux_001_src23_endofpacket),   //          .endofpacket
		.src24_ready         (cmd_xbar_demux_001_src24_ready),         //     src24.ready
		.src24_valid         (cmd_xbar_demux_001_src24_valid),         //          .valid
		.src24_data          (cmd_xbar_demux_001_src24_data),          //          .data
		.src24_channel       (cmd_xbar_demux_001_src24_channel),       //          .channel
		.src24_startofpacket (cmd_xbar_demux_001_src24_startofpacket), //          .startofpacket
		.src24_endofpacket   (cmd_xbar_demux_001_src24_endofpacket),   //          .endofpacket
		.src25_ready         (cmd_xbar_demux_001_src25_ready),         //     src25.ready
		.src25_valid         (cmd_xbar_demux_001_src25_valid),         //          .valid
		.src25_data          (cmd_xbar_demux_001_src25_data),          //          .data
		.src25_channel       (cmd_xbar_demux_001_src25_channel),       //          .channel
		.src25_startofpacket (cmd_xbar_demux_001_src25_startofpacket), //          .startofpacket
		.src25_endofpacket   (cmd_xbar_demux_001_src25_endofpacket),   //          .endofpacket
		.src26_ready         (cmd_xbar_demux_001_src26_ready),         //     src26.ready
		.src26_valid         (cmd_xbar_demux_001_src26_valid),         //          .valid
		.src26_data          (cmd_xbar_demux_001_src26_data),          //          .data
		.src26_channel       (cmd_xbar_demux_001_src26_channel),       //          .channel
		.src26_startofpacket (cmd_xbar_demux_001_src26_startofpacket), //          .startofpacket
		.src26_endofpacket   (cmd_xbar_demux_001_src26_endofpacket),   //          .endofpacket
		.src27_ready         (cmd_xbar_demux_001_src27_ready),         //     src27.ready
		.src27_valid         (cmd_xbar_demux_001_src27_valid),         //          .valid
		.src27_data          (cmd_xbar_demux_001_src27_data),          //          .data
		.src27_channel       (cmd_xbar_demux_001_src27_channel),       //          .channel
		.src27_startofpacket (cmd_xbar_demux_001_src27_startofpacket), //          .startofpacket
		.src27_endofpacket   (cmd_xbar_demux_001_src27_endofpacket),   //          .endofpacket
		.src28_ready         (cmd_xbar_demux_001_src28_ready),         //     src28.ready
		.src28_valid         (cmd_xbar_demux_001_src28_valid),         //          .valid
		.src28_data          (cmd_xbar_demux_001_src28_data),          //          .data
		.src28_channel       (cmd_xbar_demux_001_src28_channel),       //          .channel
		.src28_startofpacket (cmd_xbar_demux_001_src28_startofpacket), //          .startofpacket
		.src28_endofpacket   (cmd_xbar_demux_001_src28_endofpacket),   //          .endofpacket
		.src29_ready         (cmd_xbar_demux_001_src29_ready),         //     src29.ready
		.src29_valid         (cmd_xbar_demux_001_src29_valid),         //          .valid
		.src29_data          (cmd_xbar_demux_001_src29_data),          //          .data
		.src29_channel       (cmd_xbar_demux_001_src29_channel),       //          .channel
		.src29_startofpacket (cmd_xbar_demux_001_src29_startofpacket), //          .startofpacket
		.src29_endofpacket   (cmd_xbar_demux_001_src29_endofpacket),   //          .endofpacket
		.src30_ready         (cmd_xbar_demux_001_src30_ready),         //     src30.ready
		.src30_valid         (cmd_xbar_demux_001_src30_valid),         //          .valid
		.src30_data          (cmd_xbar_demux_001_src30_data),          //          .data
		.src30_channel       (cmd_xbar_demux_001_src30_channel),       //          .channel
		.src30_startofpacket (cmd_xbar_demux_001_src30_startofpacket), //          .startofpacket
		.src30_endofpacket   (cmd_xbar_demux_001_src30_endofpacket),   //          .endofpacket
		.src31_ready         (cmd_xbar_demux_001_src31_ready),         //     src31.ready
		.src31_valid         (cmd_xbar_demux_001_src31_valid),         //          .valid
		.src31_data          (cmd_xbar_demux_001_src31_data),          //          .data
		.src31_channel       (cmd_xbar_demux_001_src31_channel),       //          .channel
		.src31_startofpacket (cmd_xbar_demux_001_src31_startofpacket), //          .startofpacket
		.src31_endofpacket   (cmd_xbar_demux_001_src31_endofpacket),   //          .endofpacket
		.src32_ready         (cmd_xbar_demux_001_src32_ready),         //     src32.ready
		.src32_valid         (cmd_xbar_demux_001_src32_valid),         //          .valid
		.src32_data          (cmd_xbar_demux_001_src32_data),          //          .data
		.src32_channel       (cmd_xbar_demux_001_src32_channel),       //          .channel
		.src32_startofpacket (cmd_xbar_demux_001_src32_startofpacket), //          .startofpacket
		.src32_endofpacket   (cmd_xbar_demux_001_src32_endofpacket),   //          .endofpacket
		.src33_ready         (cmd_xbar_demux_001_src33_ready),         //     src33.ready
		.src33_valid         (cmd_xbar_demux_001_src33_valid),         //          .valid
		.src33_data          (cmd_xbar_demux_001_src33_data),          //          .data
		.src33_channel       (cmd_xbar_demux_001_src33_channel),       //          .channel
		.src33_startofpacket (cmd_xbar_demux_001_src33_startofpacket), //          .startofpacket
		.src33_endofpacket   (cmd_xbar_demux_001_src33_endofpacket),   //          .endofpacket
		.src34_ready         (cmd_xbar_demux_001_src34_ready),         //     src34.ready
		.src34_valid         (cmd_xbar_demux_001_src34_valid),         //          .valid
		.src34_data          (cmd_xbar_demux_001_src34_data),          //          .data
		.src34_channel       (cmd_xbar_demux_001_src34_channel),       //          .channel
		.src34_startofpacket (cmd_xbar_demux_001_src34_startofpacket), //          .startofpacket
		.src34_endofpacket   (cmd_xbar_demux_001_src34_endofpacket),   //          .endofpacket
		.src35_ready         (cmd_xbar_demux_001_src35_ready),         //     src35.ready
		.src35_valid         (cmd_xbar_demux_001_src35_valid),         //          .valid
		.src35_data          (cmd_xbar_demux_001_src35_data),          //          .data
		.src35_channel       (cmd_xbar_demux_001_src35_channel),       //          .channel
		.src35_startofpacket (cmd_xbar_demux_001_src35_startofpacket), //          .startofpacket
		.src35_endofpacket   (cmd_xbar_demux_001_src35_endofpacket),   //          .endofpacket
		.src36_ready         (cmd_xbar_demux_001_src36_ready),         //     src36.ready
		.src36_valid         (cmd_xbar_demux_001_src36_valid),         //          .valid
		.src36_data          (cmd_xbar_demux_001_src36_data),          //          .data
		.src36_channel       (cmd_xbar_demux_001_src36_channel),       //          .channel
		.src36_startofpacket (cmd_xbar_demux_001_src36_startofpacket), //          .startofpacket
		.src36_endofpacket   (cmd_xbar_demux_001_src36_endofpacket),   //          .endofpacket
		.src37_ready         (cmd_xbar_demux_001_src37_ready),         //     src37.ready
		.src37_valid         (cmd_xbar_demux_001_src37_valid),         //          .valid
		.src37_data          (cmd_xbar_demux_001_src37_data),          //          .data
		.src37_channel       (cmd_xbar_demux_001_src37_channel),       //          .channel
		.src37_startofpacket (cmd_xbar_demux_001_src37_startofpacket), //          .startofpacket
		.src37_endofpacket   (cmd_xbar_demux_001_src37_endofpacket),   //          .endofpacket
		.src38_ready         (cmd_xbar_demux_001_src38_ready),         //     src38.ready
		.src38_valid         (cmd_xbar_demux_001_src38_valid),         //          .valid
		.src38_data          (cmd_xbar_demux_001_src38_data),          //          .data
		.src38_channel       (cmd_xbar_demux_001_src38_channel),       //          .channel
		.src38_startofpacket (cmd_xbar_demux_001_src38_startofpacket), //          .startofpacket
		.src38_endofpacket   (cmd_xbar_demux_001_src38_endofpacket),   //          .endofpacket
		.src39_ready         (cmd_xbar_demux_001_src39_ready),         //     src39.ready
		.src39_valid         (cmd_xbar_demux_001_src39_valid),         //          .valid
		.src39_data          (cmd_xbar_demux_001_src39_data),          //          .data
		.src39_channel       (cmd_xbar_demux_001_src39_channel),       //          .channel
		.src39_startofpacket (cmd_xbar_demux_001_src39_startofpacket), //          .startofpacket
		.src39_endofpacket   (cmd_xbar_demux_001_src39_endofpacket),   //          .endofpacket
		.src40_ready         (cmd_xbar_demux_001_src40_ready),         //     src40.ready
		.src40_valid         (cmd_xbar_demux_001_src40_valid),         //          .valid
		.src40_data          (cmd_xbar_demux_001_src40_data),          //          .data
		.src40_channel       (cmd_xbar_demux_001_src40_channel),       //          .channel
		.src40_startofpacket (cmd_xbar_demux_001_src40_startofpacket), //          .startofpacket
		.src40_endofpacket   (cmd_xbar_demux_001_src40_endofpacket),   //          .endofpacket
		.src41_ready         (cmd_xbar_demux_001_src41_ready),         //     src41.ready
		.src41_valid         (cmd_xbar_demux_001_src41_valid),         //          .valid
		.src41_data          (cmd_xbar_demux_001_src41_data),          //          .data
		.src41_channel       (cmd_xbar_demux_001_src41_channel),       //          .channel
		.src41_startofpacket (cmd_xbar_demux_001_src41_startofpacket), //          .startofpacket
		.src41_endofpacket   (cmd_xbar_demux_001_src41_endofpacket),   //          .endofpacket
		.src42_ready         (cmd_xbar_demux_001_src42_ready),         //     src42.ready
		.src42_valid         (cmd_xbar_demux_001_src42_valid),         //          .valid
		.src42_data          (cmd_xbar_demux_001_src42_data),          //          .data
		.src42_channel       (cmd_xbar_demux_001_src42_channel),       //          .channel
		.src42_startofpacket (cmd_xbar_demux_001_src42_startofpacket), //          .startofpacket
		.src42_endofpacket   (cmd_xbar_demux_001_src42_endofpacket),   //          .endofpacket
		.src43_ready         (cmd_xbar_demux_001_src43_ready),         //     src43.ready
		.src43_valid         (cmd_xbar_demux_001_src43_valid),         //          .valid
		.src43_data          (cmd_xbar_demux_001_src43_data),          //          .data
		.src43_channel       (cmd_xbar_demux_001_src43_channel),       //          .channel
		.src43_startofpacket (cmd_xbar_demux_001_src43_startofpacket), //          .startofpacket
		.src43_endofpacket   (cmd_xbar_demux_001_src43_endofpacket),   //          .endofpacket
		.src44_ready         (cmd_xbar_demux_001_src44_ready),         //     src44.ready
		.src44_valid         (cmd_xbar_demux_001_src44_valid),         //          .valid
		.src44_data          (cmd_xbar_demux_001_src44_data),          //          .data
		.src44_channel       (cmd_xbar_demux_001_src44_channel),       //          .channel
		.src44_startofpacket (cmd_xbar_demux_001_src44_startofpacket), //          .startofpacket
		.src44_endofpacket   (cmd_xbar_demux_001_src44_endofpacket),   //          .endofpacket
		.src45_ready         (cmd_xbar_demux_001_src45_ready),         //     src45.ready
		.src45_valid         (cmd_xbar_demux_001_src45_valid),         //          .valid
		.src45_data          (cmd_xbar_demux_001_src45_data),          //          .data
		.src45_channel       (cmd_xbar_demux_001_src45_channel),       //          .channel
		.src45_startofpacket (cmd_xbar_demux_001_src45_startofpacket), //          .startofpacket
		.src45_endofpacket   (cmd_xbar_demux_001_src45_endofpacket),   //          .endofpacket
		.src46_ready         (cmd_xbar_demux_001_src46_ready),         //     src46.ready
		.src46_valid         (cmd_xbar_demux_001_src46_valid),         //          .valid
		.src46_data          (cmd_xbar_demux_001_src46_data),          //          .data
		.src46_channel       (cmd_xbar_demux_001_src46_channel),       //          .channel
		.src46_startofpacket (cmd_xbar_demux_001_src46_startofpacket), //          .startofpacket
		.src46_endofpacket   (cmd_xbar_demux_001_src46_endofpacket),   //          .endofpacket
		.src47_ready         (cmd_xbar_demux_001_src47_ready),         //     src47.ready
		.src47_valid         (cmd_xbar_demux_001_src47_valid),         //          .valid
		.src47_data          (cmd_xbar_demux_001_src47_data),          //          .data
		.src47_channel       (cmd_xbar_demux_001_src47_channel),       //          .channel
		.src47_startofpacket (cmd_xbar_demux_001_src47_startofpacket), //          .startofpacket
		.src47_endofpacket   (cmd_xbar_demux_001_src47_endofpacket),   //          .endofpacket
		.src48_ready         (cmd_xbar_demux_001_src48_ready),         //     src48.ready
		.src48_valid         (cmd_xbar_demux_001_src48_valid),         //          .valid
		.src48_data          (cmd_xbar_demux_001_src48_data),          //          .data
		.src48_channel       (cmd_xbar_demux_001_src48_channel),       //          .channel
		.src48_startofpacket (cmd_xbar_demux_001_src48_startofpacket), //          .startofpacket
		.src48_endofpacket   (cmd_xbar_demux_001_src48_endofpacket),   //          .endofpacket
		.src49_ready         (cmd_xbar_demux_001_src49_ready),         //     src49.ready
		.src49_valid         (cmd_xbar_demux_001_src49_valid),         //          .valid
		.src49_data          (cmd_xbar_demux_001_src49_data),          //          .data
		.src49_channel       (cmd_xbar_demux_001_src49_channel),       //          .channel
		.src49_startofpacket (cmd_xbar_demux_001_src49_startofpacket), //          .startofpacket
		.src49_endofpacket   (cmd_xbar_demux_001_src49_endofpacket),   //          .endofpacket
		.src50_ready         (cmd_xbar_demux_001_src50_ready),         //     src50.ready
		.src50_valid         (cmd_xbar_demux_001_src50_valid),         //          .valid
		.src50_data          (cmd_xbar_demux_001_src50_data),          //          .data
		.src50_channel       (cmd_xbar_demux_001_src50_channel),       //          .channel
		.src50_startofpacket (cmd_xbar_demux_001_src50_startofpacket), //          .startofpacket
		.src50_endofpacket   (cmd_xbar_demux_001_src50_endofpacket),   //          .endofpacket
		.src51_ready         (cmd_xbar_demux_001_src51_ready),         //     src51.ready
		.src51_valid         (cmd_xbar_demux_001_src51_valid),         //          .valid
		.src51_data          (cmd_xbar_demux_001_src51_data),          //          .data
		.src51_channel       (cmd_xbar_demux_001_src51_channel),       //          .channel
		.src51_startofpacket (cmd_xbar_demux_001_src51_startofpacket), //          .startofpacket
		.src51_endofpacket   (cmd_xbar_demux_001_src51_endofpacket),   //          .endofpacket
		.src52_ready         (cmd_xbar_demux_001_src52_ready),         //     src52.ready
		.src52_valid         (cmd_xbar_demux_001_src52_valid),         //          .valid
		.src52_data          (cmd_xbar_demux_001_src52_data),          //          .data
		.src52_channel       (cmd_xbar_demux_001_src52_channel),       //          .channel
		.src52_startofpacket (cmd_xbar_demux_001_src52_startofpacket), //          .startofpacket
		.src52_endofpacket   (cmd_xbar_demux_001_src52_endofpacket),   //          .endofpacket
		.src53_ready         (cmd_xbar_demux_001_src53_ready),         //     src53.ready
		.src53_valid         (cmd_xbar_demux_001_src53_valid),         //          .valid
		.src53_data          (cmd_xbar_demux_001_src53_data),          //          .data
		.src53_channel       (cmd_xbar_demux_001_src53_channel),       //          .channel
		.src53_startofpacket (cmd_xbar_demux_001_src53_startofpacket), //          .startofpacket
		.src53_endofpacket   (cmd_xbar_demux_001_src53_endofpacket),   //          .endofpacket
		.src54_ready         (cmd_xbar_demux_001_src54_ready),         //     src54.ready
		.src54_valid         (cmd_xbar_demux_001_src54_valid),         //          .valid
		.src54_data          (cmd_xbar_demux_001_src54_data),          //          .data
		.src54_channel       (cmd_xbar_demux_001_src54_channel),       //          .channel
		.src54_startofpacket (cmd_xbar_demux_001_src54_startofpacket), //          .startofpacket
		.src54_endofpacket   (cmd_xbar_demux_001_src54_endofpacket),   //          .endofpacket
		.src55_ready         (cmd_xbar_demux_001_src55_ready),         //     src55.ready
		.src55_valid         (cmd_xbar_demux_001_src55_valid),         //          .valid
		.src55_data          (cmd_xbar_demux_001_src55_data),          //          .data
		.src55_channel       (cmd_xbar_demux_001_src55_channel),       //          .channel
		.src55_startofpacket (cmd_xbar_demux_001_src55_startofpacket), //          .startofpacket
		.src55_endofpacket   (cmd_xbar_demux_001_src55_endofpacket),   //          .endofpacket
		.src56_ready         (cmd_xbar_demux_001_src56_ready),         //     src56.ready
		.src56_valid         (cmd_xbar_demux_001_src56_valid),         //          .valid
		.src56_data          (cmd_xbar_demux_001_src56_data),          //          .data
		.src56_channel       (cmd_xbar_demux_001_src56_channel),       //          .channel
		.src56_startofpacket (cmd_xbar_demux_001_src56_startofpacket), //          .startofpacket
		.src56_endofpacket   (cmd_xbar_demux_001_src56_endofpacket),   //          .endofpacket
		.src57_ready         (cmd_xbar_demux_001_src57_ready),         //     src57.ready
		.src57_valid         (cmd_xbar_demux_001_src57_valid),         //          .valid
		.src57_data          (cmd_xbar_demux_001_src57_data),          //          .data
		.src57_channel       (cmd_xbar_demux_001_src57_channel),       //          .channel
		.src57_startofpacket (cmd_xbar_demux_001_src57_startofpacket), //          .startofpacket
		.src57_endofpacket   (cmd_xbar_demux_001_src57_endofpacket),   //          .endofpacket
		.src58_ready         (cmd_xbar_demux_001_src58_ready),         //     src58.ready
		.src58_valid         (cmd_xbar_demux_001_src58_valid),         //          .valid
		.src58_data          (cmd_xbar_demux_001_src58_data),          //          .data
		.src58_channel       (cmd_xbar_demux_001_src58_channel),       //          .channel
		.src58_startofpacket (cmd_xbar_demux_001_src58_startofpacket), //          .startofpacket
		.src58_endofpacket   (cmd_xbar_demux_001_src58_endofpacket),   //          .endofpacket
		.src59_ready         (cmd_xbar_demux_001_src59_ready),         //     src59.ready
		.src59_valid         (cmd_xbar_demux_001_src59_valid),         //          .valid
		.src59_data          (cmd_xbar_demux_001_src59_data),          //          .data
		.src59_channel       (cmd_xbar_demux_001_src59_channel),       //          .channel
		.src59_startofpacket (cmd_xbar_demux_001_src59_startofpacket), //          .startofpacket
		.src59_endofpacket   (cmd_xbar_demux_001_src59_endofpacket),   //          .endofpacket
		.src60_ready         (cmd_xbar_demux_001_src60_ready),         //     src60.ready
		.src60_valid         (cmd_xbar_demux_001_src60_valid),         //          .valid
		.src60_data          (cmd_xbar_demux_001_src60_data),          //          .data
		.src60_channel       (cmd_xbar_demux_001_src60_channel),       //          .channel
		.src60_startofpacket (cmd_xbar_demux_001_src60_startofpacket), //          .startofpacket
		.src60_endofpacket   (cmd_xbar_demux_001_src60_endofpacket),   //          .endofpacket
		.src61_ready         (cmd_xbar_demux_001_src61_ready),         //     src61.ready
		.src61_valid         (cmd_xbar_demux_001_src61_valid),         //          .valid
		.src61_data          (cmd_xbar_demux_001_src61_data),          //          .data
		.src61_channel       (cmd_xbar_demux_001_src61_channel),       //          .channel
		.src61_startofpacket (cmd_xbar_demux_001_src61_startofpacket), //          .startofpacket
		.src61_endofpacket   (cmd_xbar_demux_001_src61_endofpacket),   //          .endofpacket
		.src62_ready         (cmd_xbar_demux_001_src62_ready),         //     src62.ready
		.src62_valid         (cmd_xbar_demux_001_src62_valid),         //          .valid
		.src62_data          (cmd_xbar_demux_001_src62_data),          //          .data
		.src62_channel       (cmd_xbar_demux_001_src62_channel),       //          .channel
		.src62_startofpacket (cmd_xbar_demux_001_src62_startofpacket), //          .startofpacket
		.src62_endofpacket   (cmd_xbar_demux_001_src62_endofpacket),   //          .endofpacket
		.src63_ready         (cmd_xbar_demux_001_src63_ready),         //     src63.ready
		.src63_valid         (cmd_xbar_demux_001_src63_valid),         //          .valid
		.src63_data          (cmd_xbar_demux_001_src63_data),          //          .data
		.src63_channel       (cmd_xbar_demux_001_src63_channel),       //          .channel
		.src63_startofpacket (cmd_xbar_demux_001_src63_startofpacket), //          .startofpacket
		.src63_endofpacket   (cmd_xbar_demux_001_src63_endofpacket),   //          .endofpacket
		.src64_ready         (cmd_xbar_demux_001_src64_ready),         //     src64.ready
		.src64_valid         (cmd_xbar_demux_001_src64_valid),         //          .valid
		.src64_data          (cmd_xbar_demux_001_src64_data),          //          .data
		.src64_channel       (cmd_xbar_demux_001_src64_channel),       //          .channel
		.src64_startofpacket (cmd_xbar_demux_001_src64_startofpacket), //          .startofpacket
		.src64_endofpacket   (cmd_xbar_demux_001_src64_endofpacket),   //          .endofpacket
		.src65_ready         (cmd_xbar_demux_001_src65_ready),         //     src65.ready
		.src65_valid         (cmd_xbar_demux_001_src65_valid),         //          .valid
		.src65_data          (cmd_xbar_demux_001_src65_data),          //          .data
		.src65_channel       (cmd_xbar_demux_001_src65_channel),       //          .channel
		.src65_startofpacket (cmd_xbar_demux_001_src65_startofpacket), //          .startofpacket
		.src65_endofpacket   (cmd_xbar_demux_001_src65_endofpacket),   //          .endofpacket
		.src66_ready         (cmd_xbar_demux_001_src66_ready),         //     src66.ready
		.src66_valid         (cmd_xbar_demux_001_src66_valid),         //          .valid
		.src66_data          (cmd_xbar_demux_001_src66_data),          //          .data
		.src66_channel       (cmd_xbar_demux_001_src66_channel),       //          .channel
		.src66_startofpacket (cmd_xbar_demux_001_src66_startofpacket), //          .startofpacket
		.src66_endofpacket   (cmd_xbar_demux_001_src66_endofpacket),   //          .endofpacket
		.src67_ready         (cmd_xbar_demux_001_src67_ready),         //     src67.ready
		.src67_valid         (cmd_xbar_demux_001_src67_valid),         //          .valid
		.src67_data          (cmd_xbar_demux_001_src67_data),          //          .data
		.src67_channel       (cmd_xbar_demux_001_src67_channel),       //          .channel
		.src67_startofpacket (cmd_xbar_demux_001_src67_startofpacket), //          .startofpacket
		.src67_endofpacket   (cmd_xbar_demux_001_src67_endofpacket),   //          .endofpacket
		.src68_ready         (cmd_xbar_demux_001_src68_ready),         //     src68.ready
		.src68_valid         (cmd_xbar_demux_001_src68_valid),         //          .valid
		.src68_data          (cmd_xbar_demux_001_src68_data),          //          .data
		.src68_channel       (cmd_xbar_demux_001_src68_channel),       //          .channel
		.src68_startofpacket (cmd_xbar_demux_001_src68_startofpacket), //          .startofpacket
		.src68_endofpacket   (cmd_xbar_demux_001_src68_endofpacket),   //          .endofpacket
		.src69_ready         (cmd_xbar_demux_001_src69_ready),         //     src69.ready
		.src69_valid         (cmd_xbar_demux_001_src69_valid),         //          .valid
		.src69_data          (cmd_xbar_demux_001_src69_data),          //          .data
		.src69_channel       (cmd_xbar_demux_001_src69_channel),       //          .channel
		.src69_startofpacket (cmd_xbar_demux_001_src69_startofpacket), //          .startofpacket
		.src69_endofpacket   (cmd_xbar_demux_001_src69_endofpacket),   //          .endofpacket
		.src70_ready         (cmd_xbar_demux_001_src70_ready),         //     src70.ready
		.src70_valid         (cmd_xbar_demux_001_src70_valid),         //          .valid
		.src70_data          (cmd_xbar_demux_001_src70_data),          //          .data
		.src70_channel       (cmd_xbar_demux_001_src70_channel),       //          .channel
		.src70_startofpacket (cmd_xbar_demux_001_src70_startofpacket), //          .startofpacket
		.src70_endofpacket   (cmd_xbar_demux_001_src70_endofpacket),   //          .endofpacket
		.src71_ready         (cmd_xbar_demux_001_src71_ready),         //     src71.ready
		.src71_valid         (cmd_xbar_demux_001_src71_valid),         //          .valid
		.src71_data          (cmd_xbar_demux_001_src71_data),          //          .data
		.src71_channel       (cmd_xbar_demux_001_src71_channel),       //          .channel
		.src71_startofpacket (cmd_xbar_demux_001_src71_startofpacket), //          .startofpacket
		.src71_endofpacket   (cmd_xbar_demux_001_src71_endofpacket),   //          .endofpacket
		.src72_ready         (cmd_xbar_demux_001_src72_ready),         //     src72.ready
		.src72_valid         (cmd_xbar_demux_001_src72_valid),         //          .valid
		.src72_data          (cmd_xbar_demux_001_src72_data),          //          .data
		.src72_channel       (cmd_xbar_demux_001_src72_channel),       //          .channel
		.src72_startofpacket (cmd_xbar_demux_001_src72_startofpacket), //          .startofpacket
		.src72_endofpacket   (cmd_xbar_demux_001_src72_endofpacket),   //          .endofpacket
		.src73_ready         (cmd_xbar_demux_001_src73_ready),         //     src73.ready
		.src73_valid         (cmd_xbar_demux_001_src73_valid),         //          .valid
		.src73_data          (cmd_xbar_demux_001_src73_data),          //          .data
		.src73_channel       (cmd_xbar_demux_001_src73_channel),       //          .channel
		.src73_startofpacket (cmd_xbar_demux_001_src73_startofpacket), //          .startofpacket
		.src73_endofpacket   (cmd_xbar_demux_001_src73_endofpacket),   //          .endofpacket
		.src74_ready         (cmd_xbar_demux_001_src74_ready),         //     src74.ready
		.src74_valid         (cmd_xbar_demux_001_src74_valid),         //          .valid
		.src74_data          (cmd_xbar_demux_001_src74_data),          //          .data
		.src74_channel       (cmd_xbar_demux_001_src74_channel),       //          .channel
		.src74_startofpacket (cmd_xbar_demux_001_src74_startofpacket), //          .startofpacket
		.src74_endofpacket   (cmd_xbar_demux_001_src74_endofpacket),   //          .endofpacket
		.src75_ready         (cmd_xbar_demux_001_src75_ready),         //     src75.ready
		.src75_valid         (cmd_xbar_demux_001_src75_valid),         //          .valid
		.src75_data          (cmd_xbar_demux_001_src75_data),          //          .data
		.src75_channel       (cmd_xbar_demux_001_src75_channel),       //          .channel
		.src75_startofpacket (cmd_xbar_demux_001_src75_startofpacket), //          .startofpacket
		.src75_endofpacket   (cmd_xbar_demux_001_src75_endofpacket),   //          .endofpacket
		.src76_ready         (cmd_xbar_demux_001_src76_ready),         //     src76.ready
		.src76_valid         (cmd_xbar_demux_001_src76_valid),         //          .valid
		.src76_data          (cmd_xbar_demux_001_src76_data),          //          .data
		.src76_channel       (cmd_xbar_demux_001_src76_channel),       //          .channel
		.src76_startofpacket (cmd_xbar_demux_001_src76_startofpacket), //          .startofpacket
		.src76_endofpacket   (cmd_xbar_demux_001_src76_endofpacket),   //          .endofpacket
		.src77_ready         (cmd_xbar_demux_001_src77_ready),         //     src77.ready
		.src77_valid         (cmd_xbar_demux_001_src77_valid),         //          .valid
		.src77_data          (cmd_xbar_demux_001_src77_data),          //          .data
		.src77_channel       (cmd_xbar_demux_001_src77_channel),       //          .channel
		.src77_startofpacket (cmd_xbar_demux_001_src77_startofpacket), //          .startofpacket
		.src77_endofpacket   (cmd_xbar_demux_001_src77_endofpacket),   //          .endofpacket
		.src78_ready         (cmd_xbar_demux_001_src78_ready),         //     src78.ready
		.src78_valid         (cmd_xbar_demux_001_src78_valid),         //          .valid
		.src78_data          (cmd_xbar_demux_001_src78_data),          //          .data
		.src78_channel       (cmd_xbar_demux_001_src78_channel),       //          .channel
		.src78_startofpacket (cmd_xbar_demux_001_src78_startofpacket), //          .startofpacket
		.src78_endofpacket   (cmd_xbar_demux_001_src78_endofpacket),   //          .endofpacket
		.src79_ready         (cmd_xbar_demux_001_src79_ready),         //     src79.ready
		.src79_valid         (cmd_xbar_demux_001_src79_valid),         //          .valid
		.src79_data          (cmd_xbar_demux_001_src79_data),          //          .data
		.src79_channel       (cmd_xbar_demux_001_src79_channel),       //          .channel
		.src79_startofpacket (cmd_xbar_demux_001_src79_startofpacket), //          .startofpacket
		.src79_endofpacket   (cmd_xbar_demux_001_src79_endofpacket),   //          .endofpacket
		.src80_ready         (cmd_xbar_demux_001_src80_ready),         //     src80.ready
		.src80_valid         (cmd_xbar_demux_001_src80_valid),         //          .valid
		.src80_data          (cmd_xbar_demux_001_src80_data),          //          .data
		.src80_channel       (cmd_xbar_demux_001_src80_channel),       //          .channel
		.src80_startofpacket (cmd_xbar_demux_001_src80_startofpacket), //          .startofpacket
		.src80_endofpacket   (cmd_xbar_demux_001_src80_endofpacket),   //          .endofpacket
		.src81_ready         (cmd_xbar_demux_001_src81_ready),         //     src81.ready
		.src81_valid         (cmd_xbar_demux_001_src81_valid),         //          .valid
		.src81_data          (cmd_xbar_demux_001_src81_data),          //          .data
		.src81_channel       (cmd_xbar_demux_001_src81_channel),       //          .channel
		.src81_startofpacket (cmd_xbar_demux_001_src81_startofpacket), //          .startofpacket
		.src81_endofpacket   (cmd_xbar_demux_001_src81_endofpacket),   //          .endofpacket
		.src82_ready         (cmd_xbar_demux_001_src82_ready),         //     src82.ready
		.src82_valid         (cmd_xbar_demux_001_src82_valid),         //          .valid
		.src82_data          (cmd_xbar_demux_001_src82_data),          //          .data
		.src82_channel       (cmd_xbar_demux_001_src82_channel),       //          .channel
		.src82_startofpacket (cmd_xbar_demux_001_src82_startofpacket), //          .startofpacket
		.src82_endofpacket   (cmd_xbar_demux_001_src82_endofpacket),   //          .endofpacket
		.src83_ready         (cmd_xbar_demux_001_src83_ready),         //     src83.ready
		.src83_valid         (cmd_xbar_demux_001_src83_valid),         //          .valid
		.src83_data          (cmd_xbar_demux_001_src83_data),          //          .data
		.src83_channel       (cmd_xbar_demux_001_src83_channel),       //          .channel
		.src83_startofpacket (cmd_xbar_demux_001_src83_startofpacket), //          .startofpacket
		.src83_endofpacket   (cmd_xbar_demux_001_src83_endofpacket),   //          .endofpacket
		.src84_ready         (cmd_xbar_demux_001_src84_ready),         //     src84.ready
		.src84_valid         (cmd_xbar_demux_001_src84_valid),         //          .valid
		.src84_data          (cmd_xbar_demux_001_src84_data),          //          .data
		.src84_channel       (cmd_xbar_demux_001_src84_channel),       //          .channel
		.src84_startofpacket (cmd_xbar_demux_001_src84_startofpacket), //          .startofpacket
		.src84_endofpacket   (cmd_xbar_demux_001_src84_endofpacket),   //          .endofpacket
		.src85_ready         (cmd_xbar_demux_001_src85_ready),         //     src85.ready
		.src85_valid         (cmd_xbar_demux_001_src85_valid),         //          .valid
		.src85_data          (cmd_xbar_demux_001_src85_data),          //          .data
		.src85_channel       (cmd_xbar_demux_001_src85_channel),       //          .channel
		.src85_startofpacket (cmd_xbar_demux_001_src85_startofpacket), //          .startofpacket
		.src85_endofpacket   (cmd_xbar_demux_001_src85_endofpacket),   //          .endofpacket
		.src86_ready         (cmd_xbar_demux_001_src86_ready),         //     src86.ready
		.src86_valid         (cmd_xbar_demux_001_src86_valid),         //          .valid
		.src86_data          (cmd_xbar_demux_001_src86_data),          //          .data
		.src86_channel       (cmd_xbar_demux_001_src86_channel),       //          .channel
		.src86_startofpacket (cmd_xbar_demux_001_src86_startofpacket), //          .startofpacket
		.src86_endofpacket   (cmd_xbar_demux_001_src86_endofpacket),   //          .endofpacket
		.src87_ready         (cmd_xbar_demux_001_src87_ready),         //     src87.ready
		.src87_valid         (cmd_xbar_demux_001_src87_valid),         //          .valid
		.src87_data          (cmd_xbar_demux_001_src87_data),          //          .data
		.src87_channel       (cmd_xbar_demux_001_src87_channel),       //          .channel
		.src87_startofpacket (cmd_xbar_demux_001_src87_startofpacket), //          .startofpacket
		.src87_endofpacket   (cmd_xbar_demux_001_src87_endofpacket),   //          .endofpacket
		.src88_ready         (cmd_xbar_demux_001_src88_ready),         //     src88.ready
		.src88_valid         (cmd_xbar_demux_001_src88_valid),         //          .valid
		.src88_data          (cmd_xbar_demux_001_src88_data),          //          .data
		.src88_channel       (cmd_xbar_demux_001_src88_channel),       //          .channel
		.src88_startofpacket (cmd_xbar_demux_001_src88_startofpacket), //          .startofpacket
		.src88_endofpacket   (cmd_xbar_demux_001_src88_endofpacket),   //          .endofpacket
		.src89_ready         (cmd_xbar_demux_001_src89_ready),         //     src89.ready
		.src89_valid         (cmd_xbar_demux_001_src89_valid),         //          .valid
		.src89_data          (cmd_xbar_demux_001_src89_data),          //          .data
		.src89_channel       (cmd_xbar_demux_001_src89_channel),       //          .channel
		.src89_startofpacket (cmd_xbar_demux_001_src89_startofpacket), //          .startofpacket
		.src89_endofpacket   (cmd_xbar_demux_001_src89_endofpacket),   //          .endofpacket
		.src90_ready         (cmd_xbar_demux_001_src90_ready),         //     src90.ready
		.src90_valid         (cmd_xbar_demux_001_src90_valid),         //          .valid
		.src90_data          (cmd_xbar_demux_001_src90_data),          //          .data
		.src90_channel       (cmd_xbar_demux_001_src90_channel),       //          .channel
		.src90_startofpacket (cmd_xbar_demux_001_src90_startofpacket), //          .startofpacket
		.src90_endofpacket   (cmd_xbar_demux_001_src90_endofpacket),   //          .endofpacket
		.src91_ready         (cmd_xbar_demux_001_src91_ready),         //     src91.ready
		.src91_valid         (cmd_xbar_demux_001_src91_valid),         //          .valid
		.src91_data          (cmd_xbar_demux_001_src91_data),          //          .data
		.src91_channel       (cmd_xbar_demux_001_src91_channel),       //          .channel
		.src91_startofpacket (cmd_xbar_demux_001_src91_startofpacket), //          .startofpacket
		.src91_endofpacket   (cmd_xbar_demux_001_src91_endofpacket),   //          .endofpacket
		.src92_ready         (cmd_xbar_demux_001_src92_ready),         //     src92.ready
		.src92_valid         (cmd_xbar_demux_001_src92_valid),         //          .valid
		.src92_data          (cmd_xbar_demux_001_src92_data),          //          .data
		.src92_channel       (cmd_xbar_demux_001_src92_channel),       //          .channel
		.src92_startofpacket (cmd_xbar_demux_001_src92_startofpacket), //          .startofpacket
		.src92_endofpacket   (cmd_xbar_demux_001_src92_endofpacket),   //          .endofpacket
		.src93_ready         (cmd_xbar_demux_001_src93_ready),         //     src93.ready
		.src93_valid         (cmd_xbar_demux_001_src93_valid),         //          .valid
		.src93_data          (cmd_xbar_demux_001_src93_data),          //          .data
		.src93_channel       (cmd_xbar_demux_001_src93_channel),       //          .channel
		.src93_startofpacket (cmd_xbar_demux_001_src93_startofpacket), //          .startofpacket
		.src93_endofpacket   (cmd_xbar_demux_001_src93_endofpacket),   //          .endofpacket
		.src94_ready         (cmd_xbar_demux_001_src94_ready),         //     src94.ready
		.src94_valid         (cmd_xbar_demux_001_src94_valid),         //          .valid
		.src94_data          (cmd_xbar_demux_001_src94_data),          //          .data
		.src94_channel       (cmd_xbar_demux_001_src94_channel),       //          .channel
		.src94_startofpacket (cmd_xbar_demux_001_src94_startofpacket), //          .startofpacket
		.src94_endofpacket   (cmd_xbar_demux_001_src94_endofpacket),   //          .endofpacket
		.src95_ready         (cmd_xbar_demux_001_src95_ready),         //     src95.ready
		.src95_valid         (cmd_xbar_demux_001_src95_valid),         //          .valid
		.src95_data          (cmd_xbar_demux_001_src95_data),          //          .data
		.src95_channel       (cmd_xbar_demux_001_src95_channel),       //          .channel
		.src95_startofpacket (cmd_xbar_demux_001_src95_startofpacket), //          .startofpacket
		.src95_endofpacket   (cmd_xbar_demux_001_src95_endofpacket),   //          .endofpacket
		.src96_ready         (cmd_xbar_demux_001_src96_ready),         //     src96.ready
		.src96_valid         (cmd_xbar_demux_001_src96_valid),         //          .valid
		.src96_data          (cmd_xbar_demux_001_src96_data),          //          .data
		.src96_channel       (cmd_xbar_demux_001_src96_channel),       //          .channel
		.src96_startofpacket (cmd_xbar_demux_001_src96_startofpacket), //          .startofpacket
		.src96_endofpacket   (cmd_xbar_demux_001_src96_endofpacket),   //          .endofpacket
		.src97_ready         (cmd_xbar_demux_001_src97_ready),         //     src97.ready
		.src97_valid         (cmd_xbar_demux_001_src97_valid),         //          .valid
		.src97_data          (cmd_xbar_demux_001_src97_data),          //          .data
		.src97_channel       (cmd_xbar_demux_001_src97_channel),       //          .channel
		.src97_startofpacket (cmd_xbar_demux_001_src97_startofpacket), //          .startofpacket
		.src97_endofpacket   (cmd_xbar_demux_001_src97_endofpacket),   //          .endofpacket
		.src98_ready         (cmd_xbar_demux_001_src98_ready),         //     src98.ready
		.src98_valid         (cmd_xbar_demux_001_src98_valid),         //          .valid
		.src98_data          (cmd_xbar_demux_001_src98_data),          //          .data
		.src98_channel       (cmd_xbar_demux_001_src98_channel),       //          .channel
		.src98_startofpacket (cmd_xbar_demux_001_src98_startofpacket), //          .startofpacket
		.src98_endofpacket   (cmd_xbar_demux_001_src98_endofpacket)    //          .endofpacket
	);

	NIOS_SYSTEMV3_cmd_xbar_mux cmd_xbar_mux (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_src_ready),                //       src.ready
		.src_valid           (cmd_xbar_mux_src_valid),                //          .valid
		.src_data            (cmd_xbar_mux_src_data),                 //          .data
		.src_channel         (cmd_xbar_mux_src_channel),              //          .channel
		.src_startofpacket   (cmd_xbar_mux_src_startofpacket),        //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_src_endofpacket),          //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src0_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src0_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src0_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src0_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src0_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src0_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src0_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src0_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src0_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src0_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src0_endofpacket)    //          .endofpacket
	);

	NIOS_SYSTEMV3_cmd_xbar_mux cmd_xbar_mux_001 (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.src_ready           (cmd_xbar_mux_001_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_001_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_001_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_001_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_001_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_001_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src1_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src1_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src1_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src1_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src1_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src1_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src1_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src1_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src1_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src1_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src1_endofpacket)    //          .endofpacket
	);

	NIOS_SYSTEMV3_cmd_xbar_mux cmd_xbar_mux_002 (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.src_ready           (cmd_xbar_mux_002_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_002_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_002_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_002_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_002_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_002_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src2_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src2_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src2_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src2_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src2_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src2_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src2_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src2_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src2_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src2_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src2_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src2_endofpacket)    //          .endofpacket
	);

	NIOS_SYSTEMV3_rsp_xbar_demux rsp_xbar_demux (
		.clk                (clk_clk),                           //       clk.clk
		.reset              (rst_controller_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_src_ready),               //      sink.ready
		.sink_channel       (id_router_src_channel),             //          .channel
		.sink_data          (id_router_src_data),                //          .data
		.sink_startofpacket (id_router_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_src1_endofpacket)    //          .endofpacket
	);

	NIOS_SYSTEMV3_rsp_xbar_demux rsp_xbar_demux_001 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_001_src_ready),               //      sink.ready
		.sink_channel       (id_router_001_src_channel),             //          .channel
		.sink_data          (id_router_001_src_data),                //          .data
		.sink_startofpacket (id_router_001_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_001_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_001_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_001_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_001_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_001_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_001_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_001_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_001_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_001_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_001_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_001_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_001_src1_endofpacket)    //          .endofpacket
	);

	NIOS_SYSTEMV3_rsp_xbar_demux rsp_xbar_demux_002 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_002_src_ready),               //      sink.ready
		.sink_channel       (id_router_002_src_channel),             //          .channel
		.sink_data          (id_router_002_src_data),                //          .data
		.sink_startofpacket (id_router_002_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_002_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_002_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_002_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_002_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_002_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_002_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_002_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_002_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_002_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_002_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_002_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_002_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_002_src1_endofpacket)    //          .endofpacket
	);

	NIOS_SYSTEMV3_rsp_xbar_demux_003 rsp_xbar_demux_003 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_003_src_ready),               //      sink.ready
		.sink_channel       (id_router_003_src_channel),             //          .channel
		.sink_data          (id_router_003_src_data),                //          .data
		.sink_startofpacket (id_router_003_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_003_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_003_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_003_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_003_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_003_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_003_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_003_src0_endofpacket)    //          .endofpacket
	);

	NIOS_SYSTEMV3_rsp_xbar_demux_003 rsp_xbar_demux_004 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_004_src_ready),               //      sink.ready
		.sink_channel       (id_router_004_src_channel),             //          .channel
		.sink_data          (id_router_004_src_data),                //          .data
		.sink_startofpacket (id_router_004_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_004_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_004_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_004_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_004_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_004_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_004_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_004_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_004_src0_endofpacket)    //          .endofpacket
	);

	NIOS_SYSTEMV3_rsp_xbar_demux_003 rsp_xbar_demux_005 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_005_src_ready),               //      sink.ready
		.sink_channel       (id_router_005_src_channel),             //          .channel
		.sink_data          (id_router_005_src_data),                //          .data
		.sink_startofpacket (id_router_005_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_005_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_005_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_005_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_005_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_005_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_005_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_005_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_005_src0_endofpacket)    //          .endofpacket
	);

	NIOS_SYSTEMV3_rsp_xbar_demux_003 rsp_xbar_demux_006 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_006_src_ready),               //      sink.ready
		.sink_channel       (id_router_006_src_channel),             //          .channel
		.sink_data          (id_router_006_src_data),                //          .data
		.sink_startofpacket (id_router_006_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_006_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_006_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_006_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_006_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_006_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_006_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_006_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_006_src0_endofpacket)    //          .endofpacket
	);

	NIOS_SYSTEMV3_rsp_xbar_demux_003 rsp_xbar_demux_007 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_007_src_ready),               //      sink.ready
		.sink_channel       (id_router_007_src_channel),             //          .channel
		.sink_data          (id_router_007_src_data),                //          .data
		.sink_startofpacket (id_router_007_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_007_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_007_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_007_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_007_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_007_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_007_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_007_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_007_src0_endofpacket)    //          .endofpacket
	);

	NIOS_SYSTEMV3_rsp_xbar_demux_003 rsp_xbar_demux_008 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_008_src_ready),               //      sink.ready
		.sink_channel       (id_router_008_src_channel),             //          .channel
		.sink_data          (id_router_008_src_data),                //          .data
		.sink_startofpacket (id_router_008_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_008_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_008_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_008_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_008_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_008_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_008_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_008_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_008_src0_endofpacket)    //          .endofpacket
	);

	NIOS_SYSTEMV3_rsp_xbar_demux_003 rsp_xbar_demux_009 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_009_src_ready),               //      sink.ready
		.sink_channel       (id_router_009_src_channel),             //          .channel
		.sink_data          (id_router_009_src_data),                //          .data
		.sink_startofpacket (id_router_009_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_009_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_009_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_009_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_009_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_009_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_009_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_009_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_009_src0_endofpacket)    //          .endofpacket
	);

	NIOS_SYSTEMV3_rsp_xbar_demux_003 rsp_xbar_demux_010 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_010_src_ready),               //      sink.ready
		.sink_channel       (id_router_010_src_channel),             //          .channel
		.sink_data          (id_router_010_src_data),                //          .data
		.sink_startofpacket (id_router_010_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_010_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_010_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_010_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_010_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_010_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_010_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_010_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_010_src0_endofpacket)    //          .endofpacket
	);

	NIOS_SYSTEMV3_rsp_xbar_demux_003 rsp_xbar_demux_011 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_011_src_ready),               //      sink.ready
		.sink_channel       (id_router_011_src_channel),             //          .channel
		.sink_data          (id_router_011_src_data),                //          .data
		.sink_startofpacket (id_router_011_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_011_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_011_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_011_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_011_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_011_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_011_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_011_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_011_src0_endofpacket)    //          .endofpacket
	);

	NIOS_SYSTEMV3_rsp_xbar_demux_003 rsp_xbar_demux_012 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_012_src_ready),               //      sink.ready
		.sink_channel       (id_router_012_src_channel),             //          .channel
		.sink_data          (id_router_012_src_data),                //          .data
		.sink_startofpacket (id_router_012_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_012_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_012_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_012_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_012_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_012_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_012_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_012_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_012_src0_endofpacket)    //          .endofpacket
	);

	NIOS_SYSTEMV3_rsp_xbar_demux_003 rsp_xbar_demux_013 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_013_src_ready),               //      sink.ready
		.sink_channel       (id_router_013_src_channel),             //          .channel
		.sink_data          (id_router_013_src_data),                //          .data
		.sink_startofpacket (id_router_013_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_013_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_013_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_013_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_013_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_013_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_013_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_013_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_013_src0_endofpacket)    //          .endofpacket
	);

	NIOS_SYSTEMV3_rsp_xbar_demux_003 rsp_xbar_demux_014 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_014_src_ready),               //      sink.ready
		.sink_channel       (id_router_014_src_channel),             //          .channel
		.sink_data          (id_router_014_src_data),                //          .data
		.sink_startofpacket (id_router_014_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_014_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_014_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_014_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_014_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_014_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_014_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_014_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_014_src0_endofpacket)    //          .endofpacket
	);

	NIOS_SYSTEMV3_rsp_xbar_demux_003 rsp_xbar_demux_015 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_015_src_ready),               //      sink.ready
		.sink_channel       (id_router_015_src_channel),             //          .channel
		.sink_data          (id_router_015_src_data),                //          .data
		.sink_startofpacket (id_router_015_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_015_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_015_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_015_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_015_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_015_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_015_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_015_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_015_src0_endofpacket)    //          .endofpacket
	);

	NIOS_SYSTEMV3_rsp_xbar_demux_003 rsp_xbar_demux_016 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_016_src_ready),               //      sink.ready
		.sink_channel       (id_router_016_src_channel),             //          .channel
		.sink_data          (id_router_016_src_data),                //          .data
		.sink_startofpacket (id_router_016_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_016_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_016_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_016_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_016_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_016_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_016_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_016_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_016_src0_endofpacket)    //          .endofpacket
	);

	NIOS_SYSTEMV3_rsp_xbar_demux_003 rsp_xbar_demux_017 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_017_src_ready),               //      sink.ready
		.sink_channel       (id_router_017_src_channel),             //          .channel
		.sink_data          (id_router_017_src_data),                //          .data
		.sink_startofpacket (id_router_017_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_017_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_017_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_017_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_017_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_017_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_017_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_017_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_017_src0_endofpacket)    //          .endofpacket
	);

	NIOS_SYSTEMV3_rsp_xbar_demux_003 rsp_xbar_demux_018 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_018_src_ready),               //      sink.ready
		.sink_channel       (id_router_018_src_channel),             //          .channel
		.sink_data          (id_router_018_src_data),                //          .data
		.sink_startofpacket (id_router_018_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_018_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_018_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_018_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_018_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_018_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_018_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_018_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_018_src0_endofpacket)    //          .endofpacket
	);

	NIOS_SYSTEMV3_rsp_xbar_demux_003 rsp_xbar_demux_019 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_019_src_ready),               //      sink.ready
		.sink_channel       (id_router_019_src_channel),             //          .channel
		.sink_data          (id_router_019_src_data),                //          .data
		.sink_startofpacket (id_router_019_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_019_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_019_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_019_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_019_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_019_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_019_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_019_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_019_src0_endofpacket)    //          .endofpacket
	);

	NIOS_SYSTEMV3_rsp_xbar_demux_003 rsp_xbar_demux_020 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_020_src_ready),               //      sink.ready
		.sink_channel       (id_router_020_src_channel),             //          .channel
		.sink_data          (id_router_020_src_data),                //          .data
		.sink_startofpacket (id_router_020_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_020_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_020_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_020_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_020_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_020_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_020_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_020_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_020_src0_endofpacket)    //          .endofpacket
	);

	NIOS_SYSTEMV3_rsp_xbar_demux_003 rsp_xbar_demux_021 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_021_src_ready),               //      sink.ready
		.sink_channel       (id_router_021_src_channel),             //          .channel
		.sink_data          (id_router_021_src_data),                //          .data
		.sink_startofpacket (id_router_021_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_021_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_021_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_021_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_021_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_021_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_021_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_021_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_021_src0_endofpacket)    //          .endofpacket
	);

	NIOS_SYSTEMV3_rsp_xbar_demux_003 rsp_xbar_demux_022 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_022_src_ready),               //      sink.ready
		.sink_channel       (id_router_022_src_channel),             //          .channel
		.sink_data          (id_router_022_src_data),                //          .data
		.sink_startofpacket (id_router_022_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_022_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_022_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_022_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_022_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_022_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_022_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_022_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_022_src0_endofpacket)    //          .endofpacket
	);

	NIOS_SYSTEMV3_rsp_xbar_demux_003 rsp_xbar_demux_023 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_023_src_ready),               //      sink.ready
		.sink_channel       (id_router_023_src_channel),             //          .channel
		.sink_data          (id_router_023_src_data),                //          .data
		.sink_startofpacket (id_router_023_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_023_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_023_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_023_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_023_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_023_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_023_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_023_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_023_src0_endofpacket)    //          .endofpacket
	);

	NIOS_SYSTEMV3_rsp_xbar_demux_003 rsp_xbar_demux_024 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_024_src_ready),               //      sink.ready
		.sink_channel       (id_router_024_src_channel),             //          .channel
		.sink_data          (id_router_024_src_data),                //          .data
		.sink_startofpacket (id_router_024_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_024_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_024_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_024_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_024_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_024_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_024_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_024_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_024_src0_endofpacket)    //          .endofpacket
	);

	NIOS_SYSTEMV3_rsp_xbar_demux_003 rsp_xbar_demux_025 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_025_src_ready),               //      sink.ready
		.sink_channel       (id_router_025_src_channel),             //          .channel
		.sink_data          (id_router_025_src_data),                //          .data
		.sink_startofpacket (id_router_025_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_025_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_025_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_025_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_025_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_025_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_025_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_025_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_025_src0_endofpacket)    //          .endofpacket
	);

	NIOS_SYSTEMV3_rsp_xbar_demux_003 rsp_xbar_demux_026 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_026_src_ready),               //      sink.ready
		.sink_channel       (id_router_026_src_channel),             //          .channel
		.sink_data          (id_router_026_src_data),                //          .data
		.sink_startofpacket (id_router_026_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_026_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_026_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_026_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_026_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_026_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_026_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_026_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_026_src0_endofpacket)    //          .endofpacket
	);

	NIOS_SYSTEMV3_rsp_xbar_demux_003 rsp_xbar_demux_027 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_027_src_ready),               //      sink.ready
		.sink_channel       (id_router_027_src_channel),             //          .channel
		.sink_data          (id_router_027_src_data),                //          .data
		.sink_startofpacket (id_router_027_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_027_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_027_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_027_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_027_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_027_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_027_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_027_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_027_src0_endofpacket)    //          .endofpacket
	);

	NIOS_SYSTEMV3_rsp_xbar_demux_003 rsp_xbar_demux_028 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_028_src_ready),               //      sink.ready
		.sink_channel       (id_router_028_src_channel),             //          .channel
		.sink_data          (id_router_028_src_data),                //          .data
		.sink_startofpacket (id_router_028_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_028_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_028_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_028_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_028_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_028_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_028_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_028_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_028_src0_endofpacket)    //          .endofpacket
	);

	NIOS_SYSTEMV3_rsp_xbar_demux_003 rsp_xbar_demux_029 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_029_src_ready),               //      sink.ready
		.sink_channel       (id_router_029_src_channel),             //          .channel
		.sink_data          (id_router_029_src_data),                //          .data
		.sink_startofpacket (id_router_029_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_029_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_029_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_029_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_029_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_029_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_029_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_029_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_029_src0_endofpacket)    //          .endofpacket
	);

	NIOS_SYSTEMV3_rsp_xbar_demux_003 rsp_xbar_demux_030 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_030_src_ready),               //      sink.ready
		.sink_channel       (id_router_030_src_channel),             //          .channel
		.sink_data          (id_router_030_src_data),                //          .data
		.sink_startofpacket (id_router_030_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_030_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_030_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_030_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_030_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_030_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_030_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_030_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_030_src0_endofpacket)    //          .endofpacket
	);

	NIOS_SYSTEMV3_rsp_xbar_demux_003 rsp_xbar_demux_031 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_031_src_ready),               //      sink.ready
		.sink_channel       (id_router_031_src_channel),             //          .channel
		.sink_data          (id_router_031_src_data),                //          .data
		.sink_startofpacket (id_router_031_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_031_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_031_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_031_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_031_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_031_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_031_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_031_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_031_src0_endofpacket)    //          .endofpacket
	);

	NIOS_SYSTEMV3_rsp_xbar_demux_003 rsp_xbar_demux_032 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_032_src_ready),               //      sink.ready
		.sink_channel       (id_router_032_src_channel),             //          .channel
		.sink_data          (id_router_032_src_data),                //          .data
		.sink_startofpacket (id_router_032_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_032_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_032_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_032_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_032_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_032_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_032_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_032_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_032_src0_endofpacket)    //          .endofpacket
	);

	NIOS_SYSTEMV3_rsp_xbar_demux_003 rsp_xbar_demux_033 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_033_src_ready),               //      sink.ready
		.sink_channel       (id_router_033_src_channel),             //          .channel
		.sink_data          (id_router_033_src_data),                //          .data
		.sink_startofpacket (id_router_033_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_033_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_033_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_033_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_033_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_033_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_033_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_033_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_033_src0_endofpacket)    //          .endofpacket
	);

	NIOS_SYSTEMV3_rsp_xbar_demux_003 rsp_xbar_demux_034 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_034_src_ready),               //      sink.ready
		.sink_channel       (id_router_034_src_channel),             //          .channel
		.sink_data          (id_router_034_src_data),                //          .data
		.sink_startofpacket (id_router_034_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_034_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_034_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_034_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_034_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_034_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_034_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_034_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_034_src0_endofpacket)    //          .endofpacket
	);

	NIOS_SYSTEMV3_rsp_xbar_demux_003 rsp_xbar_demux_035 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_035_src_ready),               //      sink.ready
		.sink_channel       (id_router_035_src_channel),             //          .channel
		.sink_data          (id_router_035_src_data),                //          .data
		.sink_startofpacket (id_router_035_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_035_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_035_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_035_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_035_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_035_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_035_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_035_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_035_src0_endofpacket)    //          .endofpacket
	);

	NIOS_SYSTEMV3_rsp_xbar_demux_003 rsp_xbar_demux_036 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_036_src_ready),               //      sink.ready
		.sink_channel       (id_router_036_src_channel),             //          .channel
		.sink_data          (id_router_036_src_data),                //          .data
		.sink_startofpacket (id_router_036_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_036_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_036_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_036_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_036_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_036_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_036_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_036_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_036_src0_endofpacket)    //          .endofpacket
	);

	NIOS_SYSTEMV3_rsp_xbar_demux_003 rsp_xbar_demux_037 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_037_src_ready),               //      sink.ready
		.sink_channel       (id_router_037_src_channel),             //          .channel
		.sink_data          (id_router_037_src_data),                //          .data
		.sink_startofpacket (id_router_037_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_037_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_037_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_037_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_037_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_037_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_037_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_037_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_037_src0_endofpacket)    //          .endofpacket
	);

	NIOS_SYSTEMV3_rsp_xbar_demux_003 rsp_xbar_demux_038 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_038_src_ready),               //      sink.ready
		.sink_channel       (id_router_038_src_channel),             //          .channel
		.sink_data          (id_router_038_src_data),                //          .data
		.sink_startofpacket (id_router_038_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_038_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_038_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_038_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_038_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_038_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_038_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_038_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_038_src0_endofpacket)    //          .endofpacket
	);

	NIOS_SYSTEMV3_rsp_xbar_demux_003 rsp_xbar_demux_039 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_039_src_ready),               //      sink.ready
		.sink_channel       (id_router_039_src_channel),             //          .channel
		.sink_data          (id_router_039_src_data),                //          .data
		.sink_startofpacket (id_router_039_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_039_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_039_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_039_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_039_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_039_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_039_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_039_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_039_src0_endofpacket)    //          .endofpacket
	);

	NIOS_SYSTEMV3_rsp_xbar_demux_003 rsp_xbar_demux_040 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_040_src_ready),               //      sink.ready
		.sink_channel       (id_router_040_src_channel),             //          .channel
		.sink_data          (id_router_040_src_data),                //          .data
		.sink_startofpacket (id_router_040_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_040_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_040_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_040_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_040_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_040_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_040_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_040_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_040_src0_endofpacket)    //          .endofpacket
	);

	NIOS_SYSTEMV3_rsp_xbar_demux_003 rsp_xbar_demux_041 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_041_src_ready),               //      sink.ready
		.sink_channel       (id_router_041_src_channel),             //          .channel
		.sink_data          (id_router_041_src_data),                //          .data
		.sink_startofpacket (id_router_041_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_041_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_041_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_041_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_041_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_041_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_041_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_041_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_041_src0_endofpacket)    //          .endofpacket
	);

	NIOS_SYSTEMV3_rsp_xbar_demux_003 rsp_xbar_demux_042 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_042_src_ready),               //      sink.ready
		.sink_channel       (id_router_042_src_channel),             //          .channel
		.sink_data          (id_router_042_src_data),                //          .data
		.sink_startofpacket (id_router_042_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_042_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_042_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_042_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_042_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_042_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_042_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_042_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_042_src0_endofpacket)    //          .endofpacket
	);

	NIOS_SYSTEMV3_rsp_xbar_demux_003 rsp_xbar_demux_043 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_043_src_ready),               //      sink.ready
		.sink_channel       (id_router_043_src_channel),             //          .channel
		.sink_data          (id_router_043_src_data),                //          .data
		.sink_startofpacket (id_router_043_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_043_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_043_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_043_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_043_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_043_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_043_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_043_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_043_src0_endofpacket)    //          .endofpacket
	);

	NIOS_SYSTEMV3_rsp_xbar_demux_003 rsp_xbar_demux_044 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_044_src_ready),               //      sink.ready
		.sink_channel       (id_router_044_src_channel),             //          .channel
		.sink_data          (id_router_044_src_data),                //          .data
		.sink_startofpacket (id_router_044_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_044_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_044_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_044_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_044_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_044_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_044_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_044_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_044_src0_endofpacket)    //          .endofpacket
	);

	NIOS_SYSTEMV3_rsp_xbar_demux_003 rsp_xbar_demux_045 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_045_src_ready),               //      sink.ready
		.sink_channel       (id_router_045_src_channel),             //          .channel
		.sink_data          (id_router_045_src_data),                //          .data
		.sink_startofpacket (id_router_045_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_045_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_045_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_045_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_045_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_045_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_045_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_045_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_045_src0_endofpacket)    //          .endofpacket
	);

	NIOS_SYSTEMV3_rsp_xbar_demux_003 rsp_xbar_demux_046 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_046_src_ready),               //      sink.ready
		.sink_channel       (id_router_046_src_channel),             //          .channel
		.sink_data          (id_router_046_src_data),                //          .data
		.sink_startofpacket (id_router_046_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_046_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_046_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_046_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_046_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_046_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_046_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_046_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_046_src0_endofpacket)    //          .endofpacket
	);

	NIOS_SYSTEMV3_rsp_xbar_demux_003 rsp_xbar_demux_047 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_047_src_ready),               //      sink.ready
		.sink_channel       (id_router_047_src_channel),             //          .channel
		.sink_data          (id_router_047_src_data),                //          .data
		.sink_startofpacket (id_router_047_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_047_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_047_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_047_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_047_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_047_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_047_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_047_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_047_src0_endofpacket)    //          .endofpacket
	);

	NIOS_SYSTEMV3_rsp_xbar_demux_003 rsp_xbar_demux_048 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_048_src_ready),               //      sink.ready
		.sink_channel       (id_router_048_src_channel),             //          .channel
		.sink_data          (id_router_048_src_data),                //          .data
		.sink_startofpacket (id_router_048_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_048_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_048_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_048_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_048_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_048_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_048_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_048_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_048_src0_endofpacket)    //          .endofpacket
	);

	NIOS_SYSTEMV3_rsp_xbar_demux_003 rsp_xbar_demux_049 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_049_src_ready),               //      sink.ready
		.sink_channel       (id_router_049_src_channel),             //          .channel
		.sink_data          (id_router_049_src_data),                //          .data
		.sink_startofpacket (id_router_049_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_049_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_049_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_049_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_049_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_049_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_049_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_049_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_049_src0_endofpacket)    //          .endofpacket
	);

	NIOS_SYSTEMV3_rsp_xbar_demux_003 rsp_xbar_demux_050 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_050_src_ready),               //      sink.ready
		.sink_channel       (id_router_050_src_channel),             //          .channel
		.sink_data          (id_router_050_src_data),                //          .data
		.sink_startofpacket (id_router_050_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_050_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_050_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_050_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_050_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_050_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_050_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_050_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_050_src0_endofpacket)    //          .endofpacket
	);

	NIOS_SYSTEMV3_rsp_xbar_demux_003 rsp_xbar_demux_051 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_051_src_ready),               //      sink.ready
		.sink_channel       (id_router_051_src_channel),             //          .channel
		.sink_data          (id_router_051_src_data),                //          .data
		.sink_startofpacket (id_router_051_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_051_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_051_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_051_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_051_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_051_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_051_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_051_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_051_src0_endofpacket)    //          .endofpacket
	);

	NIOS_SYSTEMV3_rsp_xbar_demux_003 rsp_xbar_demux_052 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_052_src_ready),               //      sink.ready
		.sink_channel       (id_router_052_src_channel),             //          .channel
		.sink_data          (id_router_052_src_data),                //          .data
		.sink_startofpacket (id_router_052_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_052_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_052_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_052_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_052_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_052_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_052_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_052_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_052_src0_endofpacket)    //          .endofpacket
	);

	NIOS_SYSTEMV3_rsp_xbar_demux_003 rsp_xbar_demux_053 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_053_src_ready),               //      sink.ready
		.sink_channel       (id_router_053_src_channel),             //          .channel
		.sink_data          (id_router_053_src_data),                //          .data
		.sink_startofpacket (id_router_053_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_053_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_053_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_053_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_053_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_053_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_053_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_053_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_053_src0_endofpacket)    //          .endofpacket
	);

	NIOS_SYSTEMV3_rsp_xbar_demux_003 rsp_xbar_demux_054 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_054_src_ready),               //      sink.ready
		.sink_channel       (id_router_054_src_channel),             //          .channel
		.sink_data          (id_router_054_src_data),                //          .data
		.sink_startofpacket (id_router_054_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_054_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_054_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_054_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_054_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_054_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_054_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_054_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_054_src0_endofpacket)    //          .endofpacket
	);

	NIOS_SYSTEMV3_rsp_xbar_demux_003 rsp_xbar_demux_055 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_055_src_ready),               //      sink.ready
		.sink_channel       (id_router_055_src_channel),             //          .channel
		.sink_data          (id_router_055_src_data),                //          .data
		.sink_startofpacket (id_router_055_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_055_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_055_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_055_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_055_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_055_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_055_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_055_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_055_src0_endofpacket)    //          .endofpacket
	);

	NIOS_SYSTEMV3_rsp_xbar_demux_003 rsp_xbar_demux_056 (
		.clk                (clk_clk),                                //       clk.clk
		.reset              (nios_cpu_jtag_debug_module_reset_reset), // clk_reset.reset
		.sink_ready         (id_router_056_src_ready),                //      sink.ready
		.sink_channel       (id_router_056_src_channel),              //          .channel
		.sink_data          (id_router_056_src_data),                 //          .data
		.sink_startofpacket (id_router_056_src_startofpacket),        //          .startofpacket
		.sink_endofpacket   (id_router_056_src_endofpacket),          //          .endofpacket
		.sink_valid         (id_router_056_src_valid),                //          .valid
		.src0_ready         (rsp_xbar_demux_056_src0_ready),          //      src0.ready
		.src0_valid         (rsp_xbar_demux_056_src0_valid),          //          .valid
		.src0_data          (rsp_xbar_demux_056_src0_data),           //          .data
		.src0_channel       (rsp_xbar_demux_056_src0_channel),        //          .channel
		.src0_startofpacket (rsp_xbar_demux_056_src0_startofpacket),  //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_056_src0_endofpacket)     //          .endofpacket
	);

	NIOS_SYSTEMV3_rsp_xbar_demux_003 rsp_xbar_demux_057 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_057_src_ready),               //      sink.ready
		.sink_channel       (id_router_057_src_channel),             //          .channel
		.sink_data          (id_router_057_src_data),                //          .data
		.sink_startofpacket (id_router_057_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_057_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_057_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_057_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_057_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_057_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_057_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_057_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_057_src0_endofpacket)    //          .endofpacket
	);

	NIOS_SYSTEMV3_rsp_xbar_demux_003 rsp_xbar_demux_058 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_058_src_ready),               //      sink.ready
		.sink_channel       (id_router_058_src_channel),             //          .channel
		.sink_data          (id_router_058_src_data),                //          .data
		.sink_startofpacket (id_router_058_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_058_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_058_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_058_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_058_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_058_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_058_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_058_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_058_src0_endofpacket)    //          .endofpacket
	);

	NIOS_SYSTEMV3_rsp_xbar_demux_003 rsp_xbar_demux_059 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_059_src_ready),               //      sink.ready
		.sink_channel       (id_router_059_src_channel),             //          .channel
		.sink_data          (id_router_059_src_data),                //          .data
		.sink_startofpacket (id_router_059_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_059_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_059_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_059_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_059_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_059_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_059_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_059_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_059_src0_endofpacket)    //          .endofpacket
	);

	NIOS_SYSTEMV3_rsp_xbar_demux_003 rsp_xbar_demux_060 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_060_src_ready),               //      sink.ready
		.sink_channel       (id_router_060_src_channel),             //          .channel
		.sink_data          (id_router_060_src_data),                //          .data
		.sink_startofpacket (id_router_060_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_060_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_060_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_060_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_060_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_060_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_060_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_060_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_060_src0_endofpacket)    //          .endofpacket
	);

	NIOS_SYSTEMV3_rsp_xbar_demux_003 rsp_xbar_demux_061 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_061_src_ready),               //      sink.ready
		.sink_channel       (id_router_061_src_channel),             //          .channel
		.sink_data          (id_router_061_src_data),                //          .data
		.sink_startofpacket (id_router_061_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_061_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_061_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_061_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_061_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_061_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_061_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_061_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_061_src0_endofpacket)    //          .endofpacket
	);

	NIOS_SYSTEMV3_rsp_xbar_demux_003 rsp_xbar_demux_062 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_062_src_ready),               //      sink.ready
		.sink_channel       (id_router_062_src_channel),             //          .channel
		.sink_data          (id_router_062_src_data),                //          .data
		.sink_startofpacket (id_router_062_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_062_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_062_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_062_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_062_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_062_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_062_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_062_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_062_src0_endofpacket)    //          .endofpacket
	);

	NIOS_SYSTEMV3_rsp_xbar_demux_003 rsp_xbar_demux_063 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_063_src_ready),               //      sink.ready
		.sink_channel       (id_router_063_src_channel),             //          .channel
		.sink_data          (id_router_063_src_data),                //          .data
		.sink_startofpacket (id_router_063_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_063_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_063_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_063_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_063_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_063_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_063_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_063_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_063_src0_endofpacket)    //          .endofpacket
	);

	NIOS_SYSTEMV3_rsp_xbar_demux_003 rsp_xbar_demux_064 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_064_src_ready),               //      sink.ready
		.sink_channel       (id_router_064_src_channel),             //          .channel
		.sink_data          (id_router_064_src_data),                //          .data
		.sink_startofpacket (id_router_064_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_064_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_064_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_064_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_064_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_064_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_064_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_064_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_064_src0_endofpacket)    //          .endofpacket
	);

	NIOS_SYSTEMV3_rsp_xbar_demux_003 rsp_xbar_demux_065 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_065_src_ready),               //      sink.ready
		.sink_channel       (id_router_065_src_channel),             //          .channel
		.sink_data          (id_router_065_src_data),                //          .data
		.sink_startofpacket (id_router_065_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_065_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_065_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_065_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_065_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_065_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_065_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_065_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_065_src0_endofpacket)    //          .endofpacket
	);

	NIOS_SYSTEMV3_rsp_xbar_demux_003 rsp_xbar_demux_066 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_066_src_ready),               //      sink.ready
		.sink_channel       (id_router_066_src_channel),             //          .channel
		.sink_data          (id_router_066_src_data),                //          .data
		.sink_startofpacket (id_router_066_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_066_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_066_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_066_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_066_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_066_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_066_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_066_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_066_src0_endofpacket)    //          .endofpacket
	);

	NIOS_SYSTEMV3_rsp_xbar_demux_003 rsp_xbar_demux_067 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_067_src_ready),               //      sink.ready
		.sink_channel       (id_router_067_src_channel),             //          .channel
		.sink_data          (id_router_067_src_data),                //          .data
		.sink_startofpacket (id_router_067_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_067_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_067_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_067_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_067_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_067_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_067_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_067_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_067_src0_endofpacket)    //          .endofpacket
	);

	NIOS_SYSTEMV3_rsp_xbar_demux_003 rsp_xbar_demux_068 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_068_src_ready),               //      sink.ready
		.sink_channel       (id_router_068_src_channel),             //          .channel
		.sink_data          (id_router_068_src_data),                //          .data
		.sink_startofpacket (id_router_068_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_068_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_068_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_068_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_068_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_068_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_068_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_068_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_068_src0_endofpacket)    //          .endofpacket
	);

	NIOS_SYSTEMV3_rsp_xbar_demux_003 rsp_xbar_demux_069 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_069_src_ready),               //      sink.ready
		.sink_channel       (id_router_069_src_channel),             //          .channel
		.sink_data          (id_router_069_src_data),                //          .data
		.sink_startofpacket (id_router_069_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_069_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_069_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_069_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_069_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_069_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_069_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_069_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_069_src0_endofpacket)    //          .endofpacket
	);

	NIOS_SYSTEMV3_rsp_xbar_demux_003 rsp_xbar_demux_070 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_070_src_ready),               //      sink.ready
		.sink_channel       (id_router_070_src_channel),             //          .channel
		.sink_data          (id_router_070_src_data),                //          .data
		.sink_startofpacket (id_router_070_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_070_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_070_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_070_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_070_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_070_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_070_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_070_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_070_src0_endofpacket)    //          .endofpacket
	);

	NIOS_SYSTEMV3_rsp_xbar_demux_003 rsp_xbar_demux_071 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_071_src_ready),               //      sink.ready
		.sink_channel       (id_router_071_src_channel),             //          .channel
		.sink_data          (id_router_071_src_data),                //          .data
		.sink_startofpacket (id_router_071_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_071_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_071_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_071_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_071_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_071_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_071_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_071_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_071_src0_endofpacket)    //          .endofpacket
	);

	NIOS_SYSTEMV3_rsp_xbar_demux_003 rsp_xbar_demux_072 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_072_src_ready),               //      sink.ready
		.sink_channel       (id_router_072_src_channel),             //          .channel
		.sink_data          (id_router_072_src_data),                //          .data
		.sink_startofpacket (id_router_072_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_072_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_072_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_072_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_072_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_072_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_072_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_072_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_072_src0_endofpacket)    //          .endofpacket
	);

	NIOS_SYSTEMV3_rsp_xbar_demux_003 rsp_xbar_demux_073 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_073_src_ready),               //      sink.ready
		.sink_channel       (id_router_073_src_channel),             //          .channel
		.sink_data          (id_router_073_src_data),                //          .data
		.sink_startofpacket (id_router_073_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_073_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_073_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_073_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_073_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_073_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_073_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_073_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_073_src0_endofpacket)    //          .endofpacket
	);

	NIOS_SYSTEMV3_rsp_xbar_demux_003 rsp_xbar_demux_074 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_074_src_ready),               //      sink.ready
		.sink_channel       (id_router_074_src_channel),             //          .channel
		.sink_data          (id_router_074_src_data),                //          .data
		.sink_startofpacket (id_router_074_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_074_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_074_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_074_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_074_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_074_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_074_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_074_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_074_src0_endofpacket)    //          .endofpacket
	);

	NIOS_SYSTEMV3_rsp_xbar_demux_003 rsp_xbar_demux_075 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_075_src_ready),               //      sink.ready
		.sink_channel       (id_router_075_src_channel),             //          .channel
		.sink_data          (id_router_075_src_data),                //          .data
		.sink_startofpacket (id_router_075_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_075_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_075_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_075_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_075_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_075_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_075_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_075_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_075_src0_endofpacket)    //          .endofpacket
	);

	NIOS_SYSTEMV3_rsp_xbar_demux_003 rsp_xbar_demux_076 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_076_src_ready),               //      sink.ready
		.sink_channel       (id_router_076_src_channel),             //          .channel
		.sink_data          (id_router_076_src_data),                //          .data
		.sink_startofpacket (id_router_076_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_076_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_076_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_076_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_076_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_076_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_076_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_076_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_076_src0_endofpacket)    //          .endofpacket
	);

	NIOS_SYSTEMV3_rsp_xbar_demux_003 rsp_xbar_demux_077 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_077_src_ready),               //      sink.ready
		.sink_channel       (id_router_077_src_channel),             //          .channel
		.sink_data          (id_router_077_src_data),                //          .data
		.sink_startofpacket (id_router_077_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_077_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_077_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_077_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_077_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_077_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_077_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_077_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_077_src0_endofpacket)    //          .endofpacket
	);

	NIOS_SYSTEMV3_rsp_xbar_demux_003 rsp_xbar_demux_078 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_078_src_ready),               //      sink.ready
		.sink_channel       (id_router_078_src_channel),             //          .channel
		.sink_data          (id_router_078_src_data),                //          .data
		.sink_startofpacket (id_router_078_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_078_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_078_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_078_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_078_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_078_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_078_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_078_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_078_src0_endofpacket)    //          .endofpacket
	);

	NIOS_SYSTEMV3_rsp_xbar_demux_003 rsp_xbar_demux_079 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_079_src_ready),               //      sink.ready
		.sink_channel       (id_router_079_src_channel),             //          .channel
		.sink_data          (id_router_079_src_data),                //          .data
		.sink_startofpacket (id_router_079_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_079_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_079_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_079_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_079_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_079_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_079_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_079_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_079_src0_endofpacket)    //          .endofpacket
	);

	NIOS_SYSTEMV3_rsp_xbar_demux_003 rsp_xbar_demux_080 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_080_src_ready),               //      sink.ready
		.sink_channel       (id_router_080_src_channel),             //          .channel
		.sink_data          (id_router_080_src_data),                //          .data
		.sink_startofpacket (id_router_080_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_080_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_080_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_080_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_080_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_080_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_080_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_080_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_080_src0_endofpacket)    //          .endofpacket
	);

	NIOS_SYSTEMV3_rsp_xbar_demux_003 rsp_xbar_demux_081 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_081_src_ready),               //      sink.ready
		.sink_channel       (id_router_081_src_channel),             //          .channel
		.sink_data          (id_router_081_src_data),                //          .data
		.sink_startofpacket (id_router_081_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_081_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_081_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_081_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_081_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_081_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_081_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_081_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_081_src0_endofpacket)    //          .endofpacket
	);

	NIOS_SYSTEMV3_rsp_xbar_demux_003 rsp_xbar_demux_082 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_082_src_ready),               //      sink.ready
		.sink_channel       (id_router_082_src_channel),             //          .channel
		.sink_data          (id_router_082_src_data),                //          .data
		.sink_startofpacket (id_router_082_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_082_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_082_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_082_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_082_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_082_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_082_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_082_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_082_src0_endofpacket)    //          .endofpacket
	);

	NIOS_SYSTEMV3_rsp_xbar_demux_003 rsp_xbar_demux_083 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_083_src_ready),               //      sink.ready
		.sink_channel       (id_router_083_src_channel),             //          .channel
		.sink_data          (id_router_083_src_data),                //          .data
		.sink_startofpacket (id_router_083_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_083_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_083_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_083_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_083_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_083_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_083_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_083_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_083_src0_endofpacket)    //          .endofpacket
	);

	NIOS_SYSTEMV3_rsp_xbar_demux_003 rsp_xbar_demux_084 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_084_src_ready),               //      sink.ready
		.sink_channel       (id_router_084_src_channel),             //          .channel
		.sink_data          (id_router_084_src_data),                //          .data
		.sink_startofpacket (id_router_084_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_084_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_084_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_084_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_084_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_084_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_084_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_084_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_084_src0_endofpacket)    //          .endofpacket
	);

	NIOS_SYSTEMV3_rsp_xbar_demux_003 rsp_xbar_demux_085 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_085_src_ready),               //      sink.ready
		.sink_channel       (id_router_085_src_channel),             //          .channel
		.sink_data          (id_router_085_src_data),                //          .data
		.sink_startofpacket (id_router_085_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_085_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_085_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_085_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_085_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_085_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_085_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_085_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_085_src0_endofpacket)    //          .endofpacket
	);

	NIOS_SYSTEMV3_rsp_xbar_demux_003 rsp_xbar_demux_086 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_086_src_ready),               //      sink.ready
		.sink_channel       (id_router_086_src_channel),             //          .channel
		.sink_data          (id_router_086_src_data),                //          .data
		.sink_startofpacket (id_router_086_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_086_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_086_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_086_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_086_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_086_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_086_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_086_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_086_src0_endofpacket)    //          .endofpacket
	);

	NIOS_SYSTEMV3_rsp_xbar_demux_003 rsp_xbar_demux_087 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_087_src_ready),               //      sink.ready
		.sink_channel       (id_router_087_src_channel),             //          .channel
		.sink_data          (id_router_087_src_data),                //          .data
		.sink_startofpacket (id_router_087_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_087_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_087_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_087_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_087_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_087_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_087_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_087_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_087_src0_endofpacket)    //          .endofpacket
	);

	NIOS_SYSTEMV3_rsp_xbar_demux_003 rsp_xbar_demux_088 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_088_src_ready),               //      sink.ready
		.sink_channel       (id_router_088_src_channel),             //          .channel
		.sink_data          (id_router_088_src_data),                //          .data
		.sink_startofpacket (id_router_088_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_088_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_088_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_088_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_088_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_088_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_088_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_088_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_088_src0_endofpacket)    //          .endofpacket
	);

	NIOS_SYSTEMV3_rsp_xbar_demux_003 rsp_xbar_demux_089 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_089_src_ready),               //      sink.ready
		.sink_channel       (id_router_089_src_channel),             //          .channel
		.sink_data          (id_router_089_src_data),                //          .data
		.sink_startofpacket (id_router_089_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_089_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_089_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_089_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_089_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_089_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_089_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_089_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_089_src0_endofpacket)    //          .endofpacket
	);

	NIOS_SYSTEMV3_rsp_xbar_demux_003 rsp_xbar_demux_090 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_090_src_ready),               //      sink.ready
		.sink_channel       (id_router_090_src_channel),             //          .channel
		.sink_data          (id_router_090_src_data),                //          .data
		.sink_startofpacket (id_router_090_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_090_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_090_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_090_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_090_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_090_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_090_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_090_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_090_src0_endofpacket)    //          .endofpacket
	);

	NIOS_SYSTEMV3_rsp_xbar_demux_003 rsp_xbar_demux_091 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_091_src_ready),               //      sink.ready
		.sink_channel       (id_router_091_src_channel),             //          .channel
		.sink_data          (id_router_091_src_data),                //          .data
		.sink_startofpacket (id_router_091_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_091_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_091_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_091_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_091_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_091_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_091_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_091_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_091_src0_endofpacket)    //          .endofpacket
	);

	NIOS_SYSTEMV3_rsp_xbar_demux_003 rsp_xbar_demux_092 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_092_src_ready),               //      sink.ready
		.sink_channel       (id_router_092_src_channel),             //          .channel
		.sink_data          (id_router_092_src_data),                //          .data
		.sink_startofpacket (id_router_092_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_092_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_092_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_092_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_092_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_092_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_092_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_092_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_092_src0_endofpacket)    //          .endofpacket
	);

	NIOS_SYSTEMV3_rsp_xbar_demux_003 rsp_xbar_demux_093 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_093_src_ready),               //      sink.ready
		.sink_channel       (id_router_093_src_channel),             //          .channel
		.sink_data          (id_router_093_src_data),                //          .data
		.sink_startofpacket (id_router_093_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_093_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_093_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_093_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_093_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_093_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_093_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_093_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_093_src0_endofpacket)    //          .endofpacket
	);

	NIOS_SYSTEMV3_rsp_xbar_demux_003 rsp_xbar_demux_094 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_094_src_ready),               //      sink.ready
		.sink_channel       (id_router_094_src_channel),             //          .channel
		.sink_data          (id_router_094_src_data),                //          .data
		.sink_startofpacket (id_router_094_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_094_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_094_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_094_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_094_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_094_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_094_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_094_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_094_src0_endofpacket)    //          .endofpacket
	);

	NIOS_SYSTEMV3_rsp_xbar_demux_003 rsp_xbar_demux_095 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_095_src_ready),               //      sink.ready
		.sink_channel       (id_router_095_src_channel),             //          .channel
		.sink_data          (id_router_095_src_data),                //          .data
		.sink_startofpacket (id_router_095_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_095_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_095_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_095_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_095_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_095_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_095_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_095_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_095_src0_endofpacket)    //          .endofpacket
	);

	NIOS_SYSTEMV3_rsp_xbar_demux_003 rsp_xbar_demux_096 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_096_src_ready),               //      sink.ready
		.sink_channel       (id_router_096_src_channel),             //          .channel
		.sink_data          (id_router_096_src_data),                //          .data
		.sink_startofpacket (id_router_096_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_096_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_096_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_096_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_096_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_096_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_096_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_096_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_096_src0_endofpacket)    //          .endofpacket
	);

	NIOS_SYSTEMV3_rsp_xbar_demux_003 rsp_xbar_demux_097 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_097_src_ready),               //      sink.ready
		.sink_channel       (id_router_097_src_channel),             //          .channel
		.sink_data          (id_router_097_src_data),                //          .data
		.sink_startofpacket (id_router_097_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_097_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_097_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_097_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_097_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_097_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_097_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_097_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_097_src0_endofpacket)    //          .endofpacket
	);

	NIOS_SYSTEMV3_rsp_xbar_demux_003 rsp_xbar_demux_098 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_098_src_ready),               //      sink.ready
		.sink_channel       (id_router_098_src_channel),             //          .channel
		.sink_data          (id_router_098_src_data),                //          .data
		.sink_startofpacket (id_router_098_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_098_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_098_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_098_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_098_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_098_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_098_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_098_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_098_src0_endofpacket)    //          .endofpacket
	);

	NIOS_SYSTEMV3_rsp_xbar_mux rsp_xbar_mux (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (rsp_xbar_mux_src_ready),                //       src.ready
		.src_valid           (rsp_xbar_mux_src_valid),                //          .valid
		.src_data            (rsp_xbar_mux_src_data),                 //          .data
		.src_channel         (rsp_xbar_mux_src_channel),              //          .channel
		.src_startofpacket   (rsp_xbar_mux_src_startofpacket),        //          .startofpacket
		.src_endofpacket     (rsp_xbar_mux_src_endofpacket),          //          .endofpacket
		.sink0_ready         (rsp_xbar_demux_src0_ready),             //     sink0.ready
		.sink0_valid         (rsp_xbar_demux_src0_valid),             //          .valid
		.sink0_channel       (rsp_xbar_demux_src0_channel),           //          .channel
		.sink0_data          (rsp_xbar_demux_src0_data),              //          .data
		.sink0_startofpacket (rsp_xbar_demux_src0_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (rsp_xbar_demux_src0_endofpacket),       //          .endofpacket
		.sink1_ready         (rsp_xbar_demux_001_src0_ready),         //     sink1.ready
		.sink1_valid         (rsp_xbar_demux_001_src0_valid),         //          .valid
		.sink1_channel       (rsp_xbar_demux_001_src0_channel),       //          .channel
		.sink1_data          (rsp_xbar_demux_001_src0_data),          //          .data
		.sink1_startofpacket (rsp_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (rsp_xbar_demux_001_src0_endofpacket),   //          .endofpacket
		.sink2_ready         (rsp_xbar_demux_002_src0_ready),         //     sink2.ready
		.sink2_valid         (rsp_xbar_demux_002_src0_valid),         //          .valid
		.sink2_channel       (rsp_xbar_demux_002_src0_channel),       //          .channel
		.sink2_data          (rsp_xbar_demux_002_src0_data),          //          .data
		.sink2_startofpacket (rsp_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.sink2_endofpacket   (rsp_xbar_demux_002_src0_endofpacket)    //          .endofpacket
	);

	NIOS_SYSTEMV3_rsp_xbar_mux_001 rsp_xbar_mux_001 (
		.clk                  (clk_clk),                               //       clk.clk
		.reset                (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready            (rsp_xbar_mux_001_src_ready),            //       src.ready
		.src_valid            (rsp_xbar_mux_001_src_valid),            //          .valid
		.src_data             (rsp_xbar_mux_001_src_data),             //          .data
		.src_channel          (rsp_xbar_mux_001_src_channel),          //          .channel
		.src_startofpacket    (rsp_xbar_mux_001_src_startofpacket),    //          .startofpacket
		.src_endofpacket      (rsp_xbar_mux_001_src_endofpacket),      //          .endofpacket
		.sink0_ready          (rsp_xbar_demux_src1_ready),             //     sink0.ready
		.sink0_valid          (rsp_xbar_demux_src1_valid),             //          .valid
		.sink0_channel        (rsp_xbar_demux_src1_channel),           //          .channel
		.sink0_data           (rsp_xbar_demux_src1_data),              //          .data
		.sink0_startofpacket  (rsp_xbar_demux_src1_startofpacket),     //          .startofpacket
		.sink0_endofpacket    (rsp_xbar_demux_src1_endofpacket),       //          .endofpacket
		.sink1_ready          (rsp_xbar_demux_001_src1_ready),         //     sink1.ready
		.sink1_valid          (rsp_xbar_demux_001_src1_valid),         //          .valid
		.sink1_channel        (rsp_xbar_demux_001_src1_channel),       //          .channel
		.sink1_data           (rsp_xbar_demux_001_src1_data),          //          .data
		.sink1_startofpacket  (rsp_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.sink1_endofpacket    (rsp_xbar_demux_001_src1_endofpacket),   //          .endofpacket
		.sink2_ready          (rsp_xbar_demux_002_src1_ready),         //     sink2.ready
		.sink2_valid          (rsp_xbar_demux_002_src1_valid),         //          .valid
		.sink2_channel        (rsp_xbar_demux_002_src1_channel),       //          .channel
		.sink2_data           (rsp_xbar_demux_002_src1_data),          //          .data
		.sink2_startofpacket  (rsp_xbar_demux_002_src1_startofpacket), //          .startofpacket
		.sink2_endofpacket    (rsp_xbar_demux_002_src1_endofpacket),   //          .endofpacket
		.sink3_ready          (rsp_xbar_demux_003_src0_ready),         //     sink3.ready
		.sink3_valid          (rsp_xbar_demux_003_src0_valid),         //          .valid
		.sink3_channel        (rsp_xbar_demux_003_src0_channel),       //          .channel
		.sink3_data           (rsp_xbar_demux_003_src0_data),          //          .data
		.sink3_startofpacket  (rsp_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.sink3_endofpacket    (rsp_xbar_demux_003_src0_endofpacket),   //          .endofpacket
		.sink4_ready          (rsp_xbar_demux_004_src0_ready),         //     sink4.ready
		.sink4_valid          (rsp_xbar_demux_004_src0_valid),         //          .valid
		.sink4_channel        (rsp_xbar_demux_004_src0_channel),       //          .channel
		.sink4_data           (rsp_xbar_demux_004_src0_data),          //          .data
		.sink4_startofpacket  (rsp_xbar_demux_004_src0_startofpacket), //          .startofpacket
		.sink4_endofpacket    (rsp_xbar_demux_004_src0_endofpacket),   //          .endofpacket
		.sink5_ready          (rsp_xbar_demux_005_src0_ready),         //     sink5.ready
		.sink5_valid          (rsp_xbar_demux_005_src0_valid),         //          .valid
		.sink5_channel        (rsp_xbar_demux_005_src0_channel),       //          .channel
		.sink5_data           (rsp_xbar_demux_005_src0_data),          //          .data
		.sink5_startofpacket  (rsp_xbar_demux_005_src0_startofpacket), //          .startofpacket
		.sink5_endofpacket    (rsp_xbar_demux_005_src0_endofpacket),   //          .endofpacket
		.sink6_ready          (rsp_xbar_demux_006_src0_ready),         //     sink6.ready
		.sink6_valid          (rsp_xbar_demux_006_src0_valid),         //          .valid
		.sink6_channel        (rsp_xbar_demux_006_src0_channel),       //          .channel
		.sink6_data           (rsp_xbar_demux_006_src0_data),          //          .data
		.sink6_startofpacket  (rsp_xbar_demux_006_src0_startofpacket), //          .startofpacket
		.sink6_endofpacket    (rsp_xbar_demux_006_src0_endofpacket),   //          .endofpacket
		.sink7_ready          (rsp_xbar_demux_007_src0_ready),         //     sink7.ready
		.sink7_valid          (rsp_xbar_demux_007_src0_valid),         //          .valid
		.sink7_channel        (rsp_xbar_demux_007_src0_channel),       //          .channel
		.sink7_data           (rsp_xbar_demux_007_src0_data),          //          .data
		.sink7_startofpacket  (rsp_xbar_demux_007_src0_startofpacket), //          .startofpacket
		.sink7_endofpacket    (rsp_xbar_demux_007_src0_endofpacket),   //          .endofpacket
		.sink8_ready          (rsp_xbar_demux_008_src0_ready),         //     sink8.ready
		.sink8_valid          (rsp_xbar_demux_008_src0_valid),         //          .valid
		.sink8_channel        (rsp_xbar_demux_008_src0_channel),       //          .channel
		.sink8_data           (rsp_xbar_demux_008_src0_data),          //          .data
		.sink8_startofpacket  (rsp_xbar_demux_008_src0_startofpacket), //          .startofpacket
		.sink8_endofpacket    (rsp_xbar_demux_008_src0_endofpacket),   //          .endofpacket
		.sink9_ready          (rsp_xbar_demux_009_src0_ready),         //     sink9.ready
		.sink9_valid          (rsp_xbar_demux_009_src0_valid),         //          .valid
		.sink9_channel        (rsp_xbar_demux_009_src0_channel),       //          .channel
		.sink9_data           (rsp_xbar_demux_009_src0_data),          //          .data
		.sink9_startofpacket  (rsp_xbar_demux_009_src0_startofpacket), //          .startofpacket
		.sink9_endofpacket    (rsp_xbar_demux_009_src0_endofpacket),   //          .endofpacket
		.sink10_ready         (rsp_xbar_demux_010_src0_ready),         //    sink10.ready
		.sink10_valid         (rsp_xbar_demux_010_src0_valid),         //          .valid
		.sink10_channel       (rsp_xbar_demux_010_src0_channel),       //          .channel
		.sink10_data          (rsp_xbar_demux_010_src0_data),          //          .data
		.sink10_startofpacket (rsp_xbar_demux_010_src0_startofpacket), //          .startofpacket
		.sink10_endofpacket   (rsp_xbar_demux_010_src0_endofpacket),   //          .endofpacket
		.sink11_ready         (rsp_xbar_demux_011_src0_ready),         //    sink11.ready
		.sink11_valid         (rsp_xbar_demux_011_src0_valid),         //          .valid
		.sink11_channel       (rsp_xbar_demux_011_src0_channel),       //          .channel
		.sink11_data          (rsp_xbar_demux_011_src0_data),          //          .data
		.sink11_startofpacket (rsp_xbar_demux_011_src0_startofpacket), //          .startofpacket
		.sink11_endofpacket   (rsp_xbar_demux_011_src0_endofpacket),   //          .endofpacket
		.sink12_ready         (rsp_xbar_demux_012_src0_ready),         //    sink12.ready
		.sink12_valid         (rsp_xbar_demux_012_src0_valid),         //          .valid
		.sink12_channel       (rsp_xbar_demux_012_src0_channel),       //          .channel
		.sink12_data          (rsp_xbar_demux_012_src0_data),          //          .data
		.sink12_startofpacket (rsp_xbar_demux_012_src0_startofpacket), //          .startofpacket
		.sink12_endofpacket   (rsp_xbar_demux_012_src0_endofpacket),   //          .endofpacket
		.sink13_ready         (rsp_xbar_demux_013_src0_ready),         //    sink13.ready
		.sink13_valid         (rsp_xbar_demux_013_src0_valid),         //          .valid
		.sink13_channel       (rsp_xbar_demux_013_src0_channel),       //          .channel
		.sink13_data          (rsp_xbar_demux_013_src0_data),          //          .data
		.sink13_startofpacket (rsp_xbar_demux_013_src0_startofpacket), //          .startofpacket
		.sink13_endofpacket   (rsp_xbar_demux_013_src0_endofpacket),   //          .endofpacket
		.sink14_ready         (rsp_xbar_demux_014_src0_ready),         //    sink14.ready
		.sink14_valid         (rsp_xbar_demux_014_src0_valid),         //          .valid
		.sink14_channel       (rsp_xbar_demux_014_src0_channel),       //          .channel
		.sink14_data          (rsp_xbar_demux_014_src0_data),          //          .data
		.sink14_startofpacket (rsp_xbar_demux_014_src0_startofpacket), //          .startofpacket
		.sink14_endofpacket   (rsp_xbar_demux_014_src0_endofpacket),   //          .endofpacket
		.sink15_ready         (rsp_xbar_demux_015_src0_ready),         //    sink15.ready
		.sink15_valid         (rsp_xbar_demux_015_src0_valid),         //          .valid
		.sink15_channel       (rsp_xbar_demux_015_src0_channel),       //          .channel
		.sink15_data          (rsp_xbar_demux_015_src0_data),          //          .data
		.sink15_startofpacket (rsp_xbar_demux_015_src0_startofpacket), //          .startofpacket
		.sink15_endofpacket   (rsp_xbar_demux_015_src0_endofpacket),   //          .endofpacket
		.sink16_ready         (rsp_xbar_demux_016_src0_ready),         //    sink16.ready
		.sink16_valid         (rsp_xbar_demux_016_src0_valid),         //          .valid
		.sink16_channel       (rsp_xbar_demux_016_src0_channel),       //          .channel
		.sink16_data          (rsp_xbar_demux_016_src0_data),          //          .data
		.sink16_startofpacket (rsp_xbar_demux_016_src0_startofpacket), //          .startofpacket
		.sink16_endofpacket   (rsp_xbar_demux_016_src0_endofpacket),   //          .endofpacket
		.sink17_ready         (rsp_xbar_demux_017_src0_ready),         //    sink17.ready
		.sink17_valid         (rsp_xbar_demux_017_src0_valid),         //          .valid
		.sink17_channel       (rsp_xbar_demux_017_src0_channel),       //          .channel
		.sink17_data          (rsp_xbar_demux_017_src0_data),          //          .data
		.sink17_startofpacket (rsp_xbar_demux_017_src0_startofpacket), //          .startofpacket
		.sink17_endofpacket   (rsp_xbar_demux_017_src0_endofpacket),   //          .endofpacket
		.sink18_ready         (rsp_xbar_demux_018_src0_ready),         //    sink18.ready
		.sink18_valid         (rsp_xbar_demux_018_src0_valid),         //          .valid
		.sink18_channel       (rsp_xbar_demux_018_src0_channel),       //          .channel
		.sink18_data          (rsp_xbar_demux_018_src0_data),          //          .data
		.sink18_startofpacket (rsp_xbar_demux_018_src0_startofpacket), //          .startofpacket
		.sink18_endofpacket   (rsp_xbar_demux_018_src0_endofpacket),   //          .endofpacket
		.sink19_ready         (rsp_xbar_demux_019_src0_ready),         //    sink19.ready
		.sink19_valid         (rsp_xbar_demux_019_src0_valid),         //          .valid
		.sink19_channel       (rsp_xbar_demux_019_src0_channel),       //          .channel
		.sink19_data          (rsp_xbar_demux_019_src0_data),          //          .data
		.sink19_startofpacket (rsp_xbar_demux_019_src0_startofpacket), //          .startofpacket
		.sink19_endofpacket   (rsp_xbar_demux_019_src0_endofpacket),   //          .endofpacket
		.sink20_ready         (rsp_xbar_demux_020_src0_ready),         //    sink20.ready
		.sink20_valid         (rsp_xbar_demux_020_src0_valid),         //          .valid
		.sink20_channel       (rsp_xbar_demux_020_src0_channel),       //          .channel
		.sink20_data          (rsp_xbar_demux_020_src0_data),          //          .data
		.sink20_startofpacket (rsp_xbar_demux_020_src0_startofpacket), //          .startofpacket
		.sink20_endofpacket   (rsp_xbar_demux_020_src0_endofpacket),   //          .endofpacket
		.sink21_ready         (rsp_xbar_demux_021_src0_ready),         //    sink21.ready
		.sink21_valid         (rsp_xbar_demux_021_src0_valid),         //          .valid
		.sink21_channel       (rsp_xbar_demux_021_src0_channel),       //          .channel
		.sink21_data          (rsp_xbar_demux_021_src0_data),          //          .data
		.sink21_startofpacket (rsp_xbar_demux_021_src0_startofpacket), //          .startofpacket
		.sink21_endofpacket   (rsp_xbar_demux_021_src0_endofpacket),   //          .endofpacket
		.sink22_ready         (rsp_xbar_demux_022_src0_ready),         //    sink22.ready
		.sink22_valid         (rsp_xbar_demux_022_src0_valid),         //          .valid
		.sink22_channel       (rsp_xbar_demux_022_src0_channel),       //          .channel
		.sink22_data          (rsp_xbar_demux_022_src0_data),          //          .data
		.sink22_startofpacket (rsp_xbar_demux_022_src0_startofpacket), //          .startofpacket
		.sink22_endofpacket   (rsp_xbar_demux_022_src0_endofpacket),   //          .endofpacket
		.sink23_ready         (rsp_xbar_demux_023_src0_ready),         //    sink23.ready
		.sink23_valid         (rsp_xbar_demux_023_src0_valid),         //          .valid
		.sink23_channel       (rsp_xbar_demux_023_src0_channel),       //          .channel
		.sink23_data          (rsp_xbar_demux_023_src0_data),          //          .data
		.sink23_startofpacket (rsp_xbar_demux_023_src0_startofpacket), //          .startofpacket
		.sink23_endofpacket   (rsp_xbar_demux_023_src0_endofpacket),   //          .endofpacket
		.sink24_ready         (rsp_xbar_demux_024_src0_ready),         //    sink24.ready
		.sink24_valid         (rsp_xbar_demux_024_src0_valid),         //          .valid
		.sink24_channel       (rsp_xbar_demux_024_src0_channel),       //          .channel
		.sink24_data          (rsp_xbar_demux_024_src0_data),          //          .data
		.sink24_startofpacket (rsp_xbar_demux_024_src0_startofpacket), //          .startofpacket
		.sink24_endofpacket   (rsp_xbar_demux_024_src0_endofpacket),   //          .endofpacket
		.sink25_ready         (rsp_xbar_demux_025_src0_ready),         //    sink25.ready
		.sink25_valid         (rsp_xbar_demux_025_src0_valid),         //          .valid
		.sink25_channel       (rsp_xbar_demux_025_src0_channel),       //          .channel
		.sink25_data          (rsp_xbar_demux_025_src0_data),          //          .data
		.sink25_startofpacket (rsp_xbar_demux_025_src0_startofpacket), //          .startofpacket
		.sink25_endofpacket   (rsp_xbar_demux_025_src0_endofpacket),   //          .endofpacket
		.sink26_ready         (rsp_xbar_demux_026_src0_ready),         //    sink26.ready
		.sink26_valid         (rsp_xbar_demux_026_src0_valid),         //          .valid
		.sink26_channel       (rsp_xbar_demux_026_src0_channel),       //          .channel
		.sink26_data          (rsp_xbar_demux_026_src0_data),          //          .data
		.sink26_startofpacket (rsp_xbar_demux_026_src0_startofpacket), //          .startofpacket
		.sink26_endofpacket   (rsp_xbar_demux_026_src0_endofpacket),   //          .endofpacket
		.sink27_ready         (rsp_xbar_demux_027_src0_ready),         //    sink27.ready
		.sink27_valid         (rsp_xbar_demux_027_src0_valid),         //          .valid
		.sink27_channel       (rsp_xbar_demux_027_src0_channel),       //          .channel
		.sink27_data          (rsp_xbar_demux_027_src0_data),          //          .data
		.sink27_startofpacket (rsp_xbar_demux_027_src0_startofpacket), //          .startofpacket
		.sink27_endofpacket   (rsp_xbar_demux_027_src0_endofpacket),   //          .endofpacket
		.sink28_ready         (rsp_xbar_demux_028_src0_ready),         //    sink28.ready
		.sink28_valid         (rsp_xbar_demux_028_src0_valid),         //          .valid
		.sink28_channel       (rsp_xbar_demux_028_src0_channel),       //          .channel
		.sink28_data          (rsp_xbar_demux_028_src0_data),          //          .data
		.sink28_startofpacket (rsp_xbar_demux_028_src0_startofpacket), //          .startofpacket
		.sink28_endofpacket   (rsp_xbar_demux_028_src0_endofpacket),   //          .endofpacket
		.sink29_ready         (rsp_xbar_demux_029_src0_ready),         //    sink29.ready
		.sink29_valid         (rsp_xbar_demux_029_src0_valid),         //          .valid
		.sink29_channel       (rsp_xbar_demux_029_src0_channel),       //          .channel
		.sink29_data          (rsp_xbar_demux_029_src0_data),          //          .data
		.sink29_startofpacket (rsp_xbar_demux_029_src0_startofpacket), //          .startofpacket
		.sink29_endofpacket   (rsp_xbar_demux_029_src0_endofpacket),   //          .endofpacket
		.sink30_ready         (rsp_xbar_demux_030_src0_ready),         //    sink30.ready
		.sink30_valid         (rsp_xbar_demux_030_src0_valid),         //          .valid
		.sink30_channel       (rsp_xbar_demux_030_src0_channel),       //          .channel
		.sink30_data          (rsp_xbar_demux_030_src0_data),          //          .data
		.sink30_startofpacket (rsp_xbar_demux_030_src0_startofpacket), //          .startofpacket
		.sink30_endofpacket   (rsp_xbar_demux_030_src0_endofpacket),   //          .endofpacket
		.sink31_ready         (rsp_xbar_demux_031_src0_ready),         //    sink31.ready
		.sink31_valid         (rsp_xbar_demux_031_src0_valid),         //          .valid
		.sink31_channel       (rsp_xbar_demux_031_src0_channel),       //          .channel
		.sink31_data          (rsp_xbar_demux_031_src0_data),          //          .data
		.sink31_startofpacket (rsp_xbar_demux_031_src0_startofpacket), //          .startofpacket
		.sink31_endofpacket   (rsp_xbar_demux_031_src0_endofpacket),   //          .endofpacket
		.sink32_ready         (rsp_xbar_demux_032_src0_ready),         //    sink32.ready
		.sink32_valid         (rsp_xbar_demux_032_src0_valid),         //          .valid
		.sink32_channel       (rsp_xbar_demux_032_src0_channel),       //          .channel
		.sink32_data          (rsp_xbar_demux_032_src0_data),          //          .data
		.sink32_startofpacket (rsp_xbar_demux_032_src0_startofpacket), //          .startofpacket
		.sink32_endofpacket   (rsp_xbar_demux_032_src0_endofpacket),   //          .endofpacket
		.sink33_ready         (rsp_xbar_demux_033_src0_ready),         //    sink33.ready
		.sink33_valid         (rsp_xbar_demux_033_src0_valid),         //          .valid
		.sink33_channel       (rsp_xbar_demux_033_src0_channel),       //          .channel
		.sink33_data          (rsp_xbar_demux_033_src0_data),          //          .data
		.sink33_startofpacket (rsp_xbar_demux_033_src0_startofpacket), //          .startofpacket
		.sink33_endofpacket   (rsp_xbar_demux_033_src0_endofpacket),   //          .endofpacket
		.sink34_ready         (rsp_xbar_demux_034_src0_ready),         //    sink34.ready
		.sink34_valid         (rsp_xbar_demux_034_src0_valid),         //          .valid
		.sink34_channel       (rsp_xbar_demux_034_src0_channel),       //          .channel
		.sink34_data          (rsp_xbar_demux_034_src0_data),          //          .data
		.sink34_startofpacket (rsp_xbar_demux_034_src0_startofpacket), //          .startofpacket
		.sink34_endofpacket   (rsp_xbar_demux_034_src0_endofpacket),   //          .endofpacket
		.sink35_ready         (rsp_xbar_demux_035_src0_ready),         //    sink35.ready
		.sink35_valid         (rsp_xbar_demux_035_src0_valid),         //          .valid
		.sink35_channel       (rsp_xbar_demux_035_src0_channel),       //          .channel
		.sink35_data          (rsp_xbar_demux_035_src0_data),          //          .data
		.sink35_startofpacket (rsp_xbar_demux_035_src0_startofpacket), //          .startofpacket
		.sink35_endofpacket   (rsp_xbar_demux_035_src0_endofpacket),   //          .endofpacket
		.sink36_ready         (rsp_xbar_demux_036_src0_ready),         //    sink36.ready
		.sink36_valid         (rsp_xbar_demux_036_src0_valid),         //          .valid
		.sink36_channel       (rsp_xbar_demux_036_src0_channel),       //          .channel
		.sink36_data          (rsp_xbar_demux_036_src0_data),          //          .data
		.sink36_startofpacket (rsp_xbar_demux_036_src0_startofpacket), //          .startofpacket
		.sink36_endofpacket   (rsp_xbar_demux_036_src0_endofpacket),   //          .endofpacket
		.sink37_ready         (rsp_xbar_demux_037_src0_ready),         //    sink37.ready
		.sink37_valid         (rsp_xbar_demux_037_src0_valid),         //          .valid
		.sink37_channel       (rsp_xbar_demux_037_src0_channel),       //          .channel
		.sink37_data          (rsp_xbar_demux_037_src0_data),          //          .data
		.sink37_startofpacket (rsp_xbar_demux_037_src0_startofpacket), //          .startofpacket
		.sink37_endofpacket   (rsp_xbar_demux_037_src0_endofpacket),   //          .endofpacket
		.sink38_ready         (rsp_xbar_demux_038_src0_ready),         //    sink38.ready
		.sink38_valid         (rsp_xbar_demux_038_src0_valid),         //          .valid
		.sink38_channel       (rsp_xbar_demux_038_src0_channel),       //          .channel
		.sink38_data          (rsp_xbar_demux_038_src0_data),          //          .data
		.sink38_startofpacket (rsp_xbar_demux_038_src0_startofpacket), //          .startofpacket
		.sink38_endofpacket   (rsp_xbar_demux_038_src0_endofpacket),   //          .endofpacket
		.sink39_ready         (rsp_xbar_demux_039_src0_ready),         //    sink39.ready
		.sink39_valid         (rsp_xbar_demux_039_src0_valid),         //          .valid
		.sink39_channel       (rsp_xbar_demux_039_src0_channel),       //          .channel
		.sink39_data          (rsp_xbar_demux_039_src0_data),          //          .data
		.sink39_startofpacket (rsp_xbar_demux_039_src0_startofpacket), //          .startofpacket
		.sink39_endofpacket   (rsp_xbar_demux_039_src0_endofpacket),   //          .endofpacket
		.sink40_ready         (rsp_xbar_demux_040_src0_ready),         //    sink40.ready
		.sink40_valid         (rsp_xbar_demux_040_src0_valid),         //          .valid
		.sink40_channel       (rsp_xbar_demux_040_src0_channel),       //          .channel
		.sink40_data          (rsp_xbar_demux_040_src0_data),          //          .data
		.sink40_startofpacket (rsp_xbar_demux_040_src0_startofpacket), //          .startofpacket
		.sink40_endofpacket   (rsp_xbar_demux_040_src0_endofpacket),   //          .endofpacket
		.sink41_ready         (rsp_xbar_demux_041_src0_ready),         //    sink41.ready
		.sink41_valid         (rsp_xbar_demux_041_src0_valid),         //          .valid
		.sink41_channel       (rsp_xbar_demux_041_src0_channel),       //          .channel
		.sink41_data          (rsp_xbar_demux_041_src0_data),          //          .data
		.sink41_startofpacket (rsp_xbar_demux_041_src0_startofpacket), //          .startofpacket
		.sink41_endofpacket   (rsp_xbar_demux_041_src0_endofpacket),   //          .endofpacket
		.sink42_ready         (rsp_xbar_demux_042_src0_ready),         //    sink42.ready
		.sink42_valid         (rsp_xbar_demux_042_src0_valid),         //          .valid
		.sink42_channel       (rsp_xbar_demux_042_src0_channel),       //          .channel
		.sink42_data          (rsp_xbar_demux_042_src0_data),          //          .data
		.sink42_startofpacket (rsp_xbar_demux_042_src0_startofpacket), //          .startofpacket
		.sink42_endofpacket   (rsp_xbar_demux_042_src0_endofpacket),   //          .endofpacket
		.sink43_ready         (rsp_xbar_demux_043_src0_ready),         //    sink43.ready
		.sink43_valid         (rsp_xbar_demux_043_src0_valid),         //          .valid
		.sink43_channel       (rsp_xbar_demux_043_src0_channel),       //          .channel
		.sink43_data          (rsp_xbar_demux_043_src0_data),          //          .data
		.sink43_startofpacket (rsp_xbar_demux_043_src0_startofpacket), //          .startofpacket
		.sink43_endofpacket   (rsp_xbar_demux_043_src0_endofpacket),   //          .endofpacket
		.sink44_ready         (rsp_xbar_demux_044_src0_ready),         //    sink44.ready
		.sink44_valid         (rsp_xbar_demux_044_src0_valid),         //          .valid
		.sink44_channel       (rsp_xbar_demux_044_src0_channel),       //          .channel
		.sink44_data          (rsp_xbar_demux_044_src0_data),          //          .data
		.sink44_startofpacket (rsp_xbar_demux_044_src0_startofpacket), //          .startofpacket
		.sink44_endofpacket   (rsp_xbar_demux_044_src0_endofpacket),   //          .endofpacket
		.sink45_ready         (rsp_xbar_demux_045_src0_ready),         //    sink45.ready
		.sink45_valid         (rsp_xbar_demux_045_src0_valid),         //          .valid
		.sink45_channel       (rsp_xbar_demux_045_src0_channel),       //          .channel
		.sink45_data          (rsp_xbar_demux_045_src0_data),          //          .data
		.sink45_startofpacket (rsp_xbar_demux_045_src0_startofpacket), //          .startofpacket
		.sink45_endofpacket   (rsp_xbar_demux_045_src0_endofpacket),   //          .endofpacket
		.sink46_ready         (rsp_xbar_demux_046_src0_ready),         //    sink46.ready
		.sink46_valid         (rsp_xbar_demux_046_src0_valid),         //          .valid
		.sink46_channel       (rsp_xbar_demux_046_src0_channel),       //          .channel
		.sink46_data          (rsp_xbar_demux_046_src0_data),          //          .data
		.sink46_startofpacket (rsp_xbar_demux_046_src0_startofpacket), //          .startofpacket
		.sink46_endofpacket   (rsp_xbar_demux_046_src0_endofpacket),   //          .endofpacket
		.sink47_ready         (rsp_xbar_demux_047_src0_ready),         //    sink47.ready
		.sink47_valid         (rsp_xbar_demux_047_src0_valid),         //          .valid
		.sink47_channel       (rsp_xbar_demux_047_src0_channel),       //          .channel
		.sink47_data          (rsp_xbar_demux_047_src0_data),          //          .data
		.sink47_startofpacket (rsp_xbar_demux_047_src0_startofpacket), //          .startofpacket
		.sink47_endofpacket   (rsp_xbar_demux_047_src0_endofpacket),   //          .endofpacket
		.sink48_ready         (rsp_xbar_demux_048_src0_ready),         //    sink48.ready
		.sink48_valid         (rsp_xbar_demux_048_src0_valid),         //          .valid
		.sink48_channel       (rsp_xbar_demux_048_src0_channel),       //          .channel
		.sink48_data          (rsp_xbar_demux_048_src0_data),          //          .data
		.sink48_startofpacket (rsp_xbar_demux_048_src0_startofpacket), //          .startofpacket
		.sink48_endofpacket   (rsp_xbar_demux_048_src0_endofpacket),   //          .endofpacket
		.sink49_ready         (rsp_xbar_demux_049_src0_ready),         //    sink49.ready
		.sink49_valid         (rsp_xbar_demux_049_src0_valid),         //          .valid
		.sink49_channel       (rsp_xbar_demux_049_src0_channel),       //          .channel
		.sink49_data          (rsp_xbar_demux_049_src0_data),          //          .data
		.sink49_startofpacket (rsp_xbar_demux_049_src0_startofpacket), //          .startofpacket
		.sink49_endofpacket   (rsp_xbar_demux_049_src0_endofpacket),   //          .endofpacket
		.sink50_ready         (rsp_xbar_demux_050_src0_ready),         //    sink50.ready
		.sink50_valid         (rsp_xbar_demux_050_src0_valid),         //          .valid
		.sink50_channel       (rsp_xbar_demux_050_src0_channel),       //          .channel
		.sink50_data          (rsp_xbar_demux_050_src0_data),          //          .data
		.sink50_startofpacket (rsp_xbar_demux_050_src0_startofpacket), //          .startofpacket
		.sink50_endofpacket   (rsp_xbar_demux_050_src0_endofpacket),   //          .endofpacket
		.sink51_ready         (rsp_xbar_demux_051_src0_ready),         //    sink51.ready
		.sink51_valid         (rsp_xbar_demux_051_src0_valid),         //          .valid
		.sink51_channel       (rsp_xbar_demux_051_src0_channel),       //          .channel
		.sink51_data          (rsp_xbar_demux_051_src0_data),          //          .data
		.sink51_startofpacket (rsp_xbar_demux_051_src0_startofpacket), //          .startofpacket
		.sink51_endofpacket   (rsp_xbar_demux_051_src0_endofpacket),   //          .endofpacket
		.sink52_ready         (rsp_xbar_demux_052_src0_ready),         //    sink52.ready
		.sink52_valid         (rsp_xbar_demux_052_src0_valid),         //          .valid
		.sink52_channel       (rsp_xbar_demux_052_src0_channel),       //          .channel
		.sink52_data          (rsp_xbar_demux_052_src0_data),          //          .data
		.sink52_startofpacket (rsp_xbar_demux_052_src0_startofpacket), //          .startofpacket
		.sink52_endofpacket   (rsp_xbar_demux_052_src0_endofpacket),   //          .endofpacket
		.sink53_ready         (rsp_xbar_demux_053_src0_ready),         //    sink53.ready
		.sink53_valid         (rsp_xbar_demux_053_src0_valid),         //          .valid
		.sink53_channel       (rsp_xbar_demux_053_src0_channel),       //          .channel
		.sink53_data          (rsp_xbar_demux_053_src0_data),          //          .data
		.sink53_startofpacket (rsp_xbar_demux_053_src0_startofpacket), //          .startofpacket
		.sink53_endofpacket   (rsp_xbar_demux_053_src0_endofpacket),   //          .endofpacket
		.sink54_ready         (rsp_xbar_demux_054_src0_ready),         //    sink54.ready
		.sink54_valid         (rsp_xbar_demux_054_src0_valid),         //          .valid
		.sink54_channel       (rsp_xbar_demux_054_src0_channel),       //          .channel
		.sink54_data          (rsp_xbar_demux_054_src0_data),          //          .data
		.sink54_startofpacket (rsp_xbar_demux_054_src0_startofpacket), //          .startofpacket
		.sink54_endofpacket   (rsp_xbar_demux_054_src0_endofpacket),   //          .endofpacket
		.sink55_ready         (rsp_xbar_demux_055_src0_ready),         //    sink55.ready
		.sink55_valid         (rsp_xbar_demux_055_src0_valid),         //          .valid
		.sink55_channel       (rsp_xbar_demux_055_src0_channel),       //          .channel
		.sink55_data          (rsp_xbar_demux_055_src0_data),          //          .data
		.sink55_startofpacket (rsp_xbar_demux_055_src0_startofpacket), //          .startofpacket
		.sink55_endofpacket   (rsp_xbar_demux_055_src0_endofpacket),   //          .endofpacket
		.sink56_ready         (rsp_xbar_demux_056_src0_ready),         //    sink56.ready
		.sink56_valid         (rsp_xbar_demux_056_src0_valid),         //          .valid
		.sink56_channel       (rsp_xbar_demux_056_src0_channel),       //          .channel
		.sink56_data          (rsp_xbar_demux_056_src0_data),          //          .data
		.sink56_startofpacket (rsp_xbar_demux_056_src0_startofpacket), //          .startofpacket
		.sink56_endofpacket   (rsp_xbar_demux_056_src0_endofpacket),   //          .endofpacket
		.sink57_ready         (rsp_xbar_demux_057_src0_ready),         //    sink57.ready
		.sink57_valid         (rsp_xbar_demux_057_src0_valid),         //          .valid
		.sink57_channel       (rsp_xbar_demux_057_src0_channel),       //          .channel
		.sink57_data          (rsp_xbar_demux_057_src0_data),          //          .data
		.sink57_startofpacket (rsp_xbar_demux_057_src0_startofpacket), //          .startofpacket
		.sink57_endofpacket   (rsp_xbar_demux_057_src0_endofpacket),   //          .endofpacket
		.sink58_ready         (rsp_xbar_demux_058_src0_ready),         //    sink58.ready
		.sink58_valid         (rsp_xbar_demux_058_src0_valid),         //          .valid
		.sink58_channel       (rsp_xbar_demux_058_src0_channel),       //          .channel
		.sink58_data          (rsp_xbar_demux_058_src0_data),          //          .data
		.sink58_startofpacket (rsp_xbar_demux_058_src0_startofpacket), //          .startofpacket
		.sink58_endofpacket   (rsp_xbar_demux_058_src0_endofpacket),   //          .endofpacket
		.sink59_ready         (rsp_xbar_demux_059_src0_ready),         //    sink59.ready
		.sink59_valid         (rsp_xbar_demux_059_src0_valid),         //          .valid
		.sink59_channel       (rsp_xbar_demux_059_src0_channel),       //          .channel
		.sink59_data          (rsp_xbar_demux_059_src0_data),          //          .data
		.sink59_startofpacket (rsp_xbar_demux_059_src0_startofpacket), //          .startofpacket
		.sink59_endofpacket   (rsp_xbar_demux_059_src0_endofpacket),   //          .endofpacket
		.sink60_ready         (rsp_xbar_demux_060_src0_ready),         //    sink60.ready
		.sink60_valid         (rsp_xbar_demux_060_src0_valid),         //          .valid
		.sink60_channel       (rsp_xbar_demux_060_src0_channel),       //          .channel
		.sink60_data          (rsp_xbar_demux_060_src0_data),          //          .data
		.sink60_startofpacket (rsp_xbar_demux_060_src0_startofpacket), //          .startofpacket
		.sink60_endofpacket   (rsp_xbar_demux_060_src0_endofpacket),   //          .endofpacket
		.sink61_ready         (rsp_xbar_demux_061_src0_ready),         //    sink61.ready
		.sink61_valid         (rsp_xbar_demux_061_src0_valid),         //          .valid
		.sink61_channel       (rsp_xbar_demux_061_src0_channel),       //          .channel
		.sink61_data          (rsp_xbar_demux_061_src0_data),          //          .data
		.sink61_startofpacket (rsp_xbar_demux_061_src0_startofpacket), //          .startofpacket
		.sink61_endofpacket   (rsp_xbar_demux_061_src0_endofpacket),   //          .endofpacket
		.sink62_ready         (rsp_xbar_demux_062_src0_ready),         //    sink62.ready
		.sink62_valid         (rsp_xbar_demux_062_src0_valid),         //          .valid
		.sink62_channel       (rsp_xbar_demux_062_src0_channel),       //          .channel
		.sink62_data          (rsp_xbar_demux_062_src0_data),          //          .data
		.sink62_startofpacket (rsp_xbar_demux_062_src0_startofpacket), //          .startofpacket
		.sink62_endofpacket   (rsp_xbar_demux_062_src0_endofpacket),   //          .endofpacket
		.sink63_ready         (rsp_xbar_demux_063_src0_ready),         //    sink63.ready
		.sink63_valid         (rsp_xbar_demux_063_src0_valid),         //          .valid
		.sink63_channel       (rsp_xbar_demux_063_src0_channel),       //          .channel
		.sink63_data          (rsp_xbar_demux_063_src0_data),          //          .data
		.sink63_startofpacket (rsp_xbar_demux_063_src0_startofpacket), //          .startofpacket
		.sink63_endofpacket   (rsp_xbar_demux_063_src0_endofpacket),   //          .endofpacket
		.sink64_ready         (rsp_xbar_demux_064_src0_ready),         //    sink64.ready
		.sink64_valid         (rsp_xbar_demux_064_src0_valid),         //          .valid
		.sink64_channel       (rsp_xbar_demux_064_src0_channel),       //          .channel
		.sink64_data          (rsp_xbar_demux_064_src0_data),          //          .data
		.sink64_startofpacket (rsp_xbar_demux_064_src0_startofpacket), //          .startofpacket
		.sink64_endofpacket   (rsp_xbar_demux_064_src0_endofpacket),   //          .endofpacket
		.sink65_ready         (rsp_xbar_demux_065_src0_ready),         //    sink65.ready
		.sink65_valid         (rsp_xbar_demux_065_src0_valid),         //          .valid
		.sink65_channel       (rsp_xbar_demux_065_src0_channel),       //          .channel
		.sink65_data          (rsp_xbar_demux_065_src0_data),          //          .data
		.sink65_startofpacket (rsp_xbar_demux_065_src0_startofpacket), //          .startofpacket
		.sink65_endofpacket   (rsp_xbar_demux_065_src0_endofpacket),   //          .endofpacket
		.sink66_ready         (rsp_xbar_demux_066_src0_ready),         //    sink66.ready
		.sink66_valid         (rsp_xbar_demux_066_src0_valid),         //          .valid
		.sink66_channel       (rsp_xbar_demux_066_src0_channel),       //          .channel
		.sink66_data          (rsp_xbar_demux_066_src0_data),          //          .data
		.sink66_startofpacket (rsp_xbar_demux_066_src0_startofpacket), //          .startofpacket
		.sink66_endofpacket   (rsp_xbar_demux_066_src0_endofpacket),   //          .endofpacket
		.sink67_ready         (rsp_xbar_demux_067_src0_ready),         //    sink67.ready
		.sink67_valid         (rsp_xbar_demux_067_src0_valid),         //          .valid
		.sink67_channel       (rsp_xbar_demux_067_src0_channel),       //          .channel
		.sink67_data          (rsp_xbar_demux_067_src0_data),          //          .data
		.sink67_startofpacket (rsp_xbar_demux_067_src0_startofpacket), //          .startofpacket
		.sink67_endofpacket   (rsp_xbar_demux_067_src0_endofpacket),   //          .endofpacket
		.sink68_ready         (rsp_xbar_demux_068_src0_ready),         //    sink68.ready
		.sink68_valid         (rsp_xbar_demux_068_src0_valid),         //          .valid
		.sink68_channel       (rsp_xbar_demux_068_src0_channel),       //          .channel
		.sink68_data          (rsp_xbar_demux_068_src0_data),          //          .data
		.sink68_startofpacket (rsp_xbar_demux_068_src0_startofpacket), //          .startofpacket
		.sink68_endofpacket   (rsp_xbar_demux_068_src0_endofpacket),   //          .endofpacket
		.sink69_ready         (rsp_xbar_demux_069_src0_ready),         //    sink69.ready
		.sink69_valid         (rsp_xbar_demux_069_src0_valid),         //          .valid
		.sink69_channel       (rsp_xbar_demux_069_src0_channel),       //          .channel
		.sink69_data          (rsp_xbar_demux_069_src0_data),          //          .data
		.sink69_startofpacket (rsp_xbar_demux_069_src0_startofpacket), //          .startofpacket
		.sink69_endofpacket   (rsp_xbar_demux_069_src0_endofpacket),   //          .endofpacket
		.sink70_ready         (rsp_xbar_demux_070_src0_ready),         //    sink70.ready
		.sink70_valid         (rsp_xbar_demux_070_src0_valid),         //          .valid
		.sink70_channel       (rsp_xbar_demux_070_src0_channel),       //          .channel
		.sink70_data          (rsp_xbar_demux_070_src0_data),          //          .data
		.sink70_startofpacket (rsp_xbar_demux_070_src0_startofpacket), //          .startofpacket
		.sink70_endofpacket   (rsp_xbar_demux_070_src0_endofpacket),   //          .endofpacket
		.sink71_ready         (rsp_xbar_demux_071_src0_ready),         //    sink71.ready
		.sink71_valid         (rsp_xbar_demux_071_src0_valid),         //          .valid
		.sink71_channel       (rsp_xbar_demux_071_src0_channel),       //          .channel
		.sink71_data          (rsp_xbar_demux_071_src0_data),          //          .data
		.sink71_startofpacket (rsp_xbar_demux_071_src0_startofpacket), //          .startofpacket
		.sink71_endofpacket   (rsp_xbar_demux_071_src0_endofpacket),   //          .endofpacket
		.sink72_ready         (rsp_xbar_demux_072_src0_ready),         //    sink72.ready
		.sink72_valid         (rsp_xbar_demux_072_src0_valid),         //          .valid
		.sink72_channel       (rsp_xbar_demux_072_src0_channel),       //          .channel
		.sink72_data          (rsp_xbar_demux_072_src0_data),          //          .data
		.sink72_startofpacket (rsp_xbar_demux_072_src0_startofpacket), //          .startofpacket
		.sink72_endofpacket   (rsp_xbar_demux_072_src0_endofpacket),   //          .endofpacket
		.sink73_ready         (rsp_xbar_demux_073_src0_ready),         //    sink73.ready
		.sink73_valid         (rsp_xbar_demux_073_src0_valid),         //          .valid
		.sink73_channel       (rsp_xbar_demux_073_src0_channel),       //          .channel
		.sink73_data          (rsp_xbar_demux_073_src0_data),          //          .data
		.sink73_startofpacket (rsp_xbar_demux_073_src0_startofpacket), //          .startofpacket
		.sink73_endofpacket   (rsp_xbar_demux_073_src0_endofpacket),   //          .endofpacket
		.sink74_ready         (rsp_xbar_demux_074_src0_ready),         //    sink74.ready
		.sink74_valid         (rsp_xbar_demux_074_src0_valid),         //          .valid
		.sink74_channel       (rsp_xbar_demux_074_src0_channel),       //          .channel
		.sink74_data          (rsp_xbar_demux_074_src0_data),          //          .data
		.sink74_startofpacket (rsp_xbar_demux_074_src0_startofpacket), //          .startofpacket
		.sink74_endofpacket   (rsp_xbar_demux_074_src0_endofpacket),   //          .endofpacket
		.sink75_ready         (rsp_xbar_demux_075_src0_ready),         //    sink75.ready
		.sink75_valid         (rsp_xbar_demux_075_src0_valid),         //          .valid
		.sink75_channel       (rsp_xbar_demux_075_src0_channel),       //          .channel
		.sink75_data          (rsp_xbar_demux_075_src0_data),          //          .data
		.sink75_startofpacket (rsp_xbar_demux_075_src0_startofpacket), //          .startofpacket
		.sink75_endofpacket   (rsp_xbar_demux_075_src0_endofpacket),   //          .endofpacket
		.sink76_ready         (rsp_xbar_demux_076_src0_ready),         //    sink76.ready
		.sink76_valid         (rsp_xbar_demux_076_src0_valid),         //          .valid
		.sink76_channel       (rsp_xbar_demux_076_src0_channel),       //          .channel
		.sink76_data          (rsp_xbar_demux_076_src0_data),          //          .data
		.sink76_startofpacket (rsp_xbar_demux_076_src0_startofpacket), //          .startofpacket
		.sink76_endofpacket   (rsp_xbar_demux_076_src0_endofpacket),   //          .endofpacket
		.sink77_ready         (rsp_xbar_demux_077_src0_ready),         //    sink77.ready
		.sink77_valid         (rsp_xbar_demux_077_src0_valid),         //          .valid
		.sink77_channel       (rsp_xbar_demux_077_src0_channel),       //          .channel
		.sink77_data          (rsp_xbar_demux_077_src0_data),          //          .data
		.sink77_startofpacket (rsp_xbar_demux_077_src0_startofpacket), //          .startofpacket
		.sink77_endofpacket   (rsp_xbar_demux_077_src0_endofpacket),   //          .endofpacket
		.sink78_ready         (rsp_xbar_demux_078_src0_ready),         //    sink78.ready
		.sink78_valid         (rsp_xbar_demux_078_src0_valid),         //          .valid
		.sink78_channel       (rsp_xbar_demux_078_src0_channel),       //          .channel
		.sink78_data          (rsp_xbar_demux_078_src0_data),          //          .data
		.sink78_startofpacket (rsp_xbar_demux_078_src0_startofpacket), //          .startofpacket
		.sink78_endofpacket   (rsp_xbar_demux_078_src0_endofpacket),   //          .endofpacket
		.sink79_ready         (rsp_xbar_demux_079_src0_ready),         //    sink79.ready
		.sink79_valid         (rsp_xbar_demux_079_src0_valid),         //          .valid
		.sink79_channel       (rsp_xbar_demux_079_src0_channel),       //          .channel
		.sink79_data          (rsp_xbar_demux_079_src0_data),          //          .data
		.sink79_startofpacket (rsp_xbar_demux_079_src0_startofpacket), //          .startofpacket
		.sink79_endofpacket   (rsp_xbar_demux_079_src0_endofpacket),   //          .endofpacket
		.sink80_ready         (rsp_xbar_demux_080_src0_ready),         //    sink80.ready
		.sink80_valid         (rsp_xbar_demux_080_src0_valid),         //          .valid
		.sink80_channel       (rsp_xbar_demux_080_src0_channel),       //          .channel
		.sink80_data          (rsp_xbar_demux_080_src0_data),          //          .data
		.sink80_startofpacket (rsp_xbar_demux_080_src0_startofpacket), //          .startofpacket
		.sink80_endofpacket   (rsp_xbar_demux_080_src0_endofpacket),   //          .endofpacket
		.sink81_ready         (rsp_xbar_demux_081_src0_ready),         //    sink81.ready
		.sink81_valid         (rsp_xbar_demux_081_src0_valid),         //          .valid
		.sink81_channel       (rsp_xbar_demux_081_src0_channel),       //          .channel
		.sink81_data          (rsp_xbar_demux_081_src0_data),          //          .data
		.sink81_startofpacket (rsp_xbar_demux_081_src0_startofpacket), //          .startofpacket
		.sink81_endofpacket   (rsp_xbar_demux_081_src0_endofpacket),   //          .endofpacket
		.sink82_ready         (rsp_xbar_demux_082_src0_ready),         //    sink82.ready
		.sink82_valid         (rsp_xbar_demux_082_src0_valid),         //          .valid
		.sink82_channel       (rsp_xbar_demux_082_src0_channel),       //          .channel
		.sink82_data          (rsp_xbar_demux_082_src0_data),          //          .data
		.sink82_startofpacket (rsp_xbar_demux_082_src0_startofpacket), //          .startofpacket
		.sink82_endofpacket   (rsp_xbar_demux_082_src0_endofpacket),   //          .endofpacket
		.sink83_ready         (rsp_xbar_demux_083_src0_ready),         //    sink83.ready
		.sink83_valid         (rsp_xbar_demux_083_src0_valid),         //          .valid
		.sink83_channel       (rsp_xbar_demux_083_src0_channel),       //          .channel
		.sink83_data          (rsp_xbar_demux_083_src0_data),          //          .data
		.sink83_startofpacket (rsp_xbar_demux_083_src0_startofpacket), //          .startofpacket
		.sink83_endofpacket   (rsp_xbar_demux_083_src0_endofpacket),   //          .endofpacket
		.sink84_ready         (rsp_xbar_demux_084_src0_ready),         //    sink84.ready
		.sink84_valid         (rsp_xbar_demux_084_src0_valid),         //          .valid
		.sink84_channel       (rsp_xbar_demux_084_src0_channel),       //          .channel
		.sink84_data          (rsp_xbar_demux_084_src0_data),          //          .data
		.sink84_startofpacket (rsp_xbar_demux_084_src0_startofpacket), //          .startofpacket
		.sink84_endofpacket   (rsp_xbar_demux_084_src0_endofpacket),   //          .endofpacket
		.sink85_ready         (rsp_xbar_demux_085_src0_ready),         //    sink85.ready
		.sink85_valid         (rsp_xbar_demux_085_src0_valid),         //          .valid
		.sink85_channel       (rsp_xbar_demux_085_src0_channel),       //          .channel
		.sink85_data          (rsp_xbar_demux_085_src0_data),          //          .data
		.sink85_startofpacket (rsp_xbar_demux_085_src0_startofpacket), //          .startofpacket
		.sink85_endofpacket   (rsp_xbar_demux_085_src0_endofpacket),   //          .endofpacket
		.sink86_ready         (rsp_xbar_demux_086_src0_ready),         //    sink86.ready
		.sink86_valid         (rsp_xbar_demux_086_src0_valid),         //          .valid
		.sink86_channel       (rsp_xbar_demux_086_src0_channel),       //          .channel
		.sink86_data          (rsp_xbar_demux_086_src0_data),          //          .data
		.sink86_startofpacket (rsp_xbar_demux_086_src0_startofpacket), //          .startofpacket
		.sink86_endofpacket   (rsp_xbar_demux_086_src0_endofpacket),   //          .endofpacket
		.sink87_ready         (rsp_xbar_demux_087_src0_ready),         //    sink87.ready
		.sink87_valid         (rsp_xbar_demux_087_src0_valid),         //          .valid
		.sink87_channel       (rsp_xbar_demux_087_src0_channel),       //          .channel
		.sink87_data          (rsp_xbar_demux_087_src0_data),          //          .data
		.sink87_startofpacket (rsp_xbar_demux_087_src0_startofpacket), //          .startofpacket
		.sink87_endofpacket   (rsp_xbar_demux_087_src0_endofpacket),   //          .endofpacket
		.sink88_ready         (rsp_xbar_demux_088_src0_ready),         //    sink88.ready
		.sink88_valid         (rsp_xbar_demux_088_src0_valid),         //          .valid
		.sink88_channel       (rsp_xbar_demux_088_src0_channel),       //          .channel
		.sink88_data          (rsp_xbar_demux_088_src0_data),          //          .data
		.sink88_startofpacket (rsp_xbar_demux_088_src0_startofpacket), //          .startofpacket
		.sink88_endofpacket   (rsp_xbar_demux_088_src0_endofpacket),   //          .endofpacket
		.sink89_ready         (rsp_xbar_demux_089_src0_ready),         //    sink89.ready
		.sink89_valid         (rsp_xbar_demux_089_src0_valid),         //          .valid
		.sink89_channel       (rsp_xbar_demux_089_src0_channel),       //          .channel
		.sink89_data          (rsp_xbar_demux_089_src0_data),          //          .data
		.sink89_startofpacket (rsp_xbar_demux_089_src0_startofpacket), //          .startofpacket
		.sink89_endofpacket   (rsp_xbar_demux_089_src0_endofpacket),   //          .endofpacket
		.sink90_ready         (rsp_xbar_demux_090_src0_ready),         //    sink90.ready
		.sink90_valid         (rsp_xbar_demux_090_src0_valid),         //          .valid
		.sink90_channel       (rsp_xbar_demux_090_src0_channel),       //          .channel
		.sink90_data          (rsp_xbar_demux_090_src0_data),          //          .data
		.sink90_startofpacket (rsp_xbar_demux_090_src0_startofpacket), //          .startofpacket
		.sink90_endofpacket   (rsp_xbar_demux_090_src0_endofpacket),   //          .endofpacket
		.sink91_ready         (rsp_xbar_demux_091_src0_ready),         //    sink91.ready
		.sink91_valid         (rsp_xbar_demux_091_src0_valid),         //          .valid
		.sink91_channel       (rsp_xbar_demux_091_src0_channel),       //          .channel
		.sink91_data          (rsp_xbar_demux_091_src0_data),          //          .data
		.sink91_startofpacket (rsp_xbar_demux_091_src0_startofpacket), //          .startofpacket
		.sink91_endofpacket   (rsp_xbar_demux_091_src0_endofpacket),   //          .endofpacket
		.sink92_ready         (rsp_xbar_demux_092_src0_ready),         //    sink92.ready
		.sink92_valid         (rsp_xbar_demux_092_src0_valid),         //          .valid
		.sink92_channel       (rsp_xbar_demux_092_src0_channel),       //          .channel
		.sink92_data          (rsp_xbar_demux_092_src0_data),          //          .data
		.sink92_startofpacket (rsp_xbar_demux_092_src0_startofpacket), //          .startofpacket
		.sink92_endofpacket   (rsp_xbar_demux_092_src0_endofpacket),   //          .endofpacket
		.sink93_ready         (rsp_xbar_demux_093_src0_ready),         //    sink93.ready
		.sink93_valid         (rsp_xbar_demux_093_src0_valid),         //          .valid
		.sink93_channel       (rsp_xbar_demux_093_src0_channel),       //          .channel
		.sink93_data          (rsp_xbar_demux_093_src0_data),          //          .data
		.sink93_startofpacket (rsp_xbar_demux_093_src0_startofpacket), //          .startofpacket
		.sink93_endofpacket   (rsp_xbar_demux_093_src0_endofpacket),   //          .endofpacket
		.sink94_ready         (rsp_xbar_demux_094_src0_ready),         //    sink94.ready
		.sink94_valid         (rsp_xbar_demux_094_src0_valid),         //          .valid
		.sink94_channel       (rsp_xbar_demux_094_src0_channel),       //          .channel
		.sink94_data          (rsp_xbar_demux_094_src0_data),          //          .data
		.sink94_startofpacket (rsp_xbar_demux_094_src0_startofpacket), //          .startofpacket
		.sink94_endofpacket   (rsp_xbar_demux_094_src0_endofpacket),   //          .endofpacket
		.sink95_ready         (rsp_xbar_demux_095_src0_ready),         //    sink95.ready
		.sink95_valid         (rsp_xbar_demux_095_src0_valid),         //          .valid
		.sink95_channel       (rsp_xbar_demux_095_src0_channel),       //          .channel
		.sink95_data          (rsp_xbar_demux_095_src0_data),          //          .data
		.sink95_startofpacket (rsp_xbar_demux_095_src0_startofpacket), //          .startofpacket
		.sink95_endofpacket   (rsp_xbar_demux_095_src0_endofpacket),   //          .endofpacket
		.sink96_ready         (rsp_xbar_demux_096_src0_ready),         //    sink96.ready
		.sink96_valid         (rsp_xbar_demux_096_src0_valid),         //          .valid
		.sink96_channel       (rsp_xbar_demux_096_src0_channel),       //          .channel
		.sink96_data          (rsp_xbar_demux_096_src0_data),          //          .data
		.sink96_startofpacket (rsp_xbar_demux_096_src0_startofpacket), //          .startofpacket
		.sink96_endofpacket   (rsp_xbar_demux_096_src0_endofpacket),   //          .endofpacket
		.sink97_ready         (rsp_xbar_demux_097_src0_ready),         //    sink97.ready
		.sink97_valid         (rsp_xbar_demux_097_src0_valid),         //          .valid
		.sink97_channel       (rsp_xbar_demux_097_src0_channel),       //          .channel
		.sink97_data          (rsp_xbar_demux_097_src0_data),          //          .data
		.sink97_startofpacket (rsp_xbar_demux_097_src0_startofpacket), //          .startofpacket
		.sink97_endofpacket   (rsp_xbar_demux_097_src0_endofpacket),   //          .endofpacket
		.sink98_ready         (rsp_xbar_demux_098_src0_ready),         //    sink98.ready
		.sink98_valid         (rsp_xbar_demux_098_src0_valid),         //          .valid
		.sink98_channel       (rsp_xbar_demux_098_src0_channel),       //          .channel
		.sink98_data          (rsp_xbar_demux_098_src0_data),          //          .data
		.sink98_startofpacket (rsp_xbar_demux_098_src0_startofpacket), //          .startofpacket
		.sink98_endofpacket   (rsp_xbar_demux_098_src0_endofpacket)    //          .endofpacket
	);

	NIOS_SYSTEMV3_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.sender_irq    (nios_cpu_d_irq_irq)              //    sender.irq
	);

endmodule
